--------------------------------------------------------------------------------
--                         Compressor_23_3_F50_uid41
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3_F50_uid41 is
    port (X1 : in  std_logic_vector(1 downto 0);
          X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3_F50_uid41 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100",
      "010" when "00011" | "00101" | "00110" | "01000" | "10000",
      "011" when "00111" | "01001" | "01010" | "01100" | "10001" | "10010" | "10100",
      "100" when "01011" | "01101" | "01110" | "10011" | "10101" | "10110" | "11000",
      "101" when "01111" | "10111" | "11001" | "11010" | "11100",
      "110" when "11011" | "11101" | "11110",
      "111" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                          Compressor_3_2_F50_uid49
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2_F50_uid49 is
    port (X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2_F50_uid49 is
signal X :  std_logic_vector(2 downto 0);
signal R0 :  std_logic_vector(1 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "00" when "000",
      "01" when "001" | "010" | "100",
      "10" when "011" | "101" | "110",
      "11" when "111",
      "--" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                         Compressor_14_3_F50_uid63
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X1 X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3_F50_uid63 is
    port (X1 : in  std_logic_vector(0 downto 0);
          X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3_F50_uid63 is
signal X :  std_logic_vector(4 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X1 & X0 ;

   with X  select  R0 <= 
      "000" when "00000",
      "001" when "00001" | "00010" | "00100" | "01000",
      "010" when "00011" | "00101" | "00110" | "01001" | "01010" | "01100" | "10000",
      "011" when "00111" | "01011" | "01101" | "01110" | "10001" | "10010" | "10100" | "11000",
      "100" when "01111" | "10011" | "10101" | "10110" | "11001" | "11010" | "11100",
      "101" when "10111" | "11011" | "11101" | "11110",
      "110" when "11111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                          Compressor_6_3_F50_uid99
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- combinatorial
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X0
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3_F50_uid99 is
    port (X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3_F50_uid99 is
signal X :  std_logic_vector(5 downto 0);
signal R0 :  std_logic_vector(2 downto 0);
begin
   X <= X0 ;

   with X  select  R0 <= 
      "000" when "000000",
      "001" when "000001" | "000010" | "000100" | "001000" | "010000" | "100000",
      "010" when "000011" | "000101" | "000110" | "001001" | "001010" | "001100" | "010001" | "010010" | "010100" | "011000" | "100001" | "100010" | "100100" | "101000" | "110000",
      "011" when "000111" | "001011" | "001101" | "001110" | "010011" | "010101" | "010110" | "011001" | "011010" | "011100" | "100011" | "100101" | "100110" | "101001" | "101010" | "101100" | "110001" | "110010" | "110100" | "111000",
      "100" when "001111" | "010111" | "011011" | "011101" | "011110" | "100111" | "101011" | "101101" | "101110" | "110011" | "110101" | "110110" | "111001" | "111010" | "111100",
      "101" when "011111" | "101111" | "110111" | "111011" | "111101" | "111110",
      "110" when "111111",
      "---" when others;
   R <= R0;
end architecture;

--------------------------------------------------------------------------------
--                      Normalizer_ZO_62_62_62_F50_uid6
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X OZb
-- Output signals: Count R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_ZO_62_62_62_F50_uid6 is
    port (clk : in std_logic;
          X : in  std_logic_vector(61 downto 0);
          OZb : in  std_logic;
          Count : out  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(61 downto 0)   );
end entity;

architecture arch of Normalizer_ZO_62_62_62_F50_uid6 is
signal level6 :  std_logic_vector(61 downto 0);
signal sozb :  std_logic;
signal count5 :  std_logic;
signal level5 :  std_logic_vector(61 downto 0);
signal count4 :  std_logic;
signal level4 :  std_logic_vector(61 downto 0);
signal count3 :  std_logic;
signal level3 :  std_logic_vector(61 downto 0);
signal count2 :  std_logic;
signal level2 :  std_logic_vector(61 downto 0);
signal count1 :  std_logic;
signal level1 :  std_logic_vector(61 downto 0);
signal count0 :  std_logic;
signal level0 :  std_logic_vector(61 downto 0);
signal sCount :  std_logic_vector(5 downto 0);
begin
   level6 <= X ;
   sozb<= OZb;
   count5<= '1' when level6(61 downto 30) = (61 downto 30=>sozb) else '0';
   level5<= level6(61 downto 0) when count5='0' else level6(29 downto 0) & (31 downto 0 => '0');

   count4<= '1' when level5(61 downto 46) = (61 downto 46=>sozb) else '0';
   level4<= level5(61 downto 0) when count4='0' else level5(45 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(61 downto 54) = (61 downto 54=>sozb) else '0';
   level3<= level4(61 downto 0) when count3='0' else level4(53 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(61 downto 58) = (61 downto 58=>sozb) else '0';
   level2<= level3(61 downto 0) when count2='0' else level3(57 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(61 downto 60) = (61 downto 60=>sozb) else '0';
   level1<= level2(61 downto 0) when count1='0' else level2(59 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(61 downto 61) = (61 downto 61=>sozb) else '0';
   level0<= level1(61 downto 0) when count0='0' else level1(60 downto 0) & (0 downto 0 => '0');

   R <= level0;
   sCount <= count5 & count4 & count3 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                       PositFastDecoder_64_2_F50_uid4
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Raul Murillo (2021)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X
-- Output signals: Sign SF Frac NZN

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity PositFastDecoder_64_2_F50_uid4 is
    port (clk : in std_logic;
          X : in  std_logic_vector(63 downto 0);
          Sign : out  std_logic;
          SF : out  std_logic_vector(8 downto 0);
          Frac : out  std_logic_vector(58 downto 0);
          NZN : out  std_logic   );
end entity;

architecture arch of PositFastDecoder_64_2_F50_uid4 is
   component Normalizer_ZO_62_62_62_F50_uid6 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(61 downto 0);
             OZb : in  std_logic;
             Count : out  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(61 downto 0)   );
   end component;

signal sgn :  std_logic;
signal pNZN :  std_logic;
signal rc :  std_logic;
signal regPosit :  std_logic_vector(61 downto 0);
signal regLength :  std_logic_vector(5 downto 0);
signal shiftedPosit :  std_logic_vector(61 downto 0);
signal k :  std_logic_vector(6 downto 0);
signal sgnVect :  std_logic_vector(1 downto 0);
signal exp :  std_logic_vector(1 downto 0);
signal pSF :  std_logic_vector(8 downto 0);
signal pFrac :  std_logic_vector(58 downto 0);
begin
--------------------------- Start of vhdl generation ---------------------------
--------------------------- Sign bit & special cases ---------------------------
   sgn <= X(63);
   pNZN <= '0' when (X(62 downto 0) = "000000000000000000000000000000000000000000000000000000000000000") else '1';
-------------- Count leading zeros/ones of regime & shift it out --------------
   rc <= X(62);
   regPosit <= X(61 downto 0);
   RegimeCounter: Normalizer_ZO_62_62_62_F50_uid6
      port map ( clk  => clk,
                 OZb => rc,
                 X => regPosit,
                 Count => regLength,
                 R => shiftedPosit);
----------------- Determine the scaling factor - regime & exp -----------------
   k <= "0" & regLength when rc /= sgn else "1" & NOT(regLength);
   sgnVect <= (others => sgn);
   exp <= shiftedPosit(60 downto 59) XOR sgnVect;
   pSF <= k & exp;
------------------------------- Extract fraction -------------------------------
   pFrac <= shiftedPosit(58 downto 0);
   Sign <= sgn;
   SF <= pSF;
   Frac <= pFrac;
   NZN <= pNZN;
---------------------------- End of vhdl generation ----------------------------
end architecture;

--------------------------------------------------------------------------------
--                      Normalizer_ZO_62_62_62_F50_uid10
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, (2007-2020)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X OZb
-- Output signals: Count R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Normalizer_ZO_62_62_62_F50_uid10 is
    port (clk : in std_logic;
          X : in  std_logic_vector(61 downto 0);
          OZb : in  std_logic;
          Count : out  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(61 downto 0)   );
end entity;

architecture arch of Normalizer_ZO_62_62_62_F50_uid10 is
signal level6 :  std_logic_vector(61 downto 0);
signal sozb :  std_logic;
signal count5 :  std_logic;
signal level5 :  std_logic_vector(61 downto 0);
signal count4 :  std_logic;
signal level4 :  std_logic_vector(61 downto 0);
signal count3 :  std_logic;
signal level3 :  std_logic_vector(61 downto 0);
signal count2 :  std_logic;
signal level2 :  std_logic_vector(61 downto 0);
signal count1 :  std_logic;
signal level1 :  std_logic_vector(61 downto 0);
signal count0 :  std_logic;
signal level0 :  std_logic_vector(61 downto 0);
signal sCount :  std_logic_vector(5 downto 0);
begin
   level6 <= X ;
   sozb<= OZb;
   count5<= '1' when level6(61 downto 30) = (61 downto 30=>sozb) else '0';
   level5<= level6(61 downto 0) when count5='0' else level6(29 downto 0) & (31 downto 0 => '0');

   count4<= '1' when level5(61 downto 46) = (61 downto 46=>sozb) else '0';
   level4<= level5(61 downto 0) when count4='0' else level5(45 downto 0) & (15 downto 0 => '0');

   count3<= '1' when level4(61 downto 54) = (61 downto 54=>sozb) else '0';
   level3<= level4(61 downto 0) when count3='0' else level4(53 downto 0) & (7 downto 0 => '0');

   count2<= '1' when level3(61 downto 58) = (61 downto 58=>sozb) else '0';
   level2<= level3(61 downto 0) when count2='0' else level3(57 downto 0) & (3 downto 0 => '0');

   count1<= '1' when level2(61 downto 60) = (61 downto 60=>sozb) else '0';
   level1<= level2(61 downto 0) when count1='0' else level2(59 downto 0) & (1 downto 0 => '0');

   count0<= '1' when level1(61 downto 61) = (61 downto 61=>sozb) else '0';
   level0<= level1(61 downto 0) when count0='0' else level1(60 downto 0) & (0 downto 0 => '0');

   R <= level0;
   sCount <= count5 & count4 & count3 & count2 & count1 & count0;
   Count <= sCount;
end architecture;

--------------------------------------------------------------------------------
--                       PositFastDecoder_64_2_F50_uid8
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Raul Murillo (2021)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X
-- Output signals: Sign SF Frac NZN

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity PositFastDecoder_64_2_F50_uid8 is
    port (clk : in std_logic;
          X : in  std_logic_vector(63 downto 0);
          Sign : out  std_logic;
          SF : out  std_logic_vector(8 downto 0);
          Frac : out  std_logic_vector(58 downto 0);
          NZN : out  std_logic   );
end entity;

architecture arch of PositFastDecoder_64_2_F50_uid8 is
   component Normalizer_ZO_62_62_62_F50_uid10 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(61 downto 0);
             OZb : in  std_logic;
             Count : out  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(61 downto 0)   );
   end component;

signal sgn :  std_logic;
signal pNZN :  std_logic;
signal rc :  std_logic;
signal regPosit :  std_logic_vector(61 downto 0);
signal regLength :  std_logic_vector(5 downto 0);
signal shiftedPosit :  std_logic_vector(61 downto 0);
signal k :  std_logic_vector(6 downto 0);
signal sgnVect :  std_logic_vector(1 downto 0);
signal exp :  std_logic_vector(1 downto 0);
signal pSF :  std_logic_vector(8 downto 0);
signal pFrac :  std_logic_vector(58 downto 0);
begin
--------------------------- Start of vhdl generation ---------------------------
--------------------------- Sign bit & special cases ---------------------------
   sgn <= X(63);
   pNZN <= '0' when (X(62 downto 0) = "000000000000000000000000000000000000000000000000000000000000000") else '1';
-------------- Count leading zeros/ones of regime & shift it out --------------
   rc <= X(62);
   regPosit <= X(61 downto 0);
   RegimeCounter: Normalizer_ZO_62_62_62_F50_uid10
      port map ( clk  => clk,
                 OZb => rc,
                 X => regPosit,
                 Count => regLength,
                 R => shiftedPosit);
----------------- Determine the scaling factor - regime & exp -----------------
   k <= "0" & regLength when rc /= sgn else "1" & NOT(regLength);
   sgnVect <= (others => sgn);
   exp <= shiftedPosit(60 downto 59) XOR sgnVect;
   pSF <= k & exp;
------------------------------- Extract fraction -------------------------------
   pFrac <= shiftedPosit(58 downto 0);
   Sign <= sgn;
   SF <= pSF;
   Frac <= pFrac;
   NZN <= pNZN;
---------------------------- End of vhdl generation ----------------------------
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_17x24_F50_uid16
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_F50_uid16 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_F50_uid16 is
signal Mint :  std_logic_vector(40 downto 0);
signal M :  std_logic_vector(40 downto 0);
signal Rtmp :  std_logic_vector(40 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(40 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_17x24_F50_uid18
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_F50_uid18 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_F50_uid18 is
signal Mint :  std_logic_vector(40 downto 0);
signal M :  std_logic_vector(40 downto 0);
signal Rtmp :  std_logic_vector(40 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(40 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_17x24_F50_uid20
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_F50_uid20 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_F50_uid20 is
signal Mint :  std_logic_vector(40 downto 0);
signal M :  std_logic_vector(40 downto 0);
signal Rtmp :  std_logic_vector(40 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(40 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_10x24_F50_uid22
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_10x24_F50_uid22 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(33 downto 0)   );
end entity;

architecture arch of DSPBlock_10x24_F50_uid22 is
signal Mint :  std_logic_vector(34 downto 0);
signal M :  std_logic_vector(33 downto 0);
signal Rtmp :  std_logic_vector(33 downto 0);
begin
   Mint <= std_logic_vector(signed(X) * signed('0' & Y)); -- multiplier
   M <= Mint(33 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_17x24_F50_uid24
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_F50_uid24 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_F50_uid24 is
signal Mint :  std_logic_vector(40 downto 0);
signal M :  std_logic_vector(40 downto 0);
signal Rtmp :  std_logic_vector(40 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(40 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_17x24_F50_uid26
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_F50_uid26 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_F50_uid26 is
signal Mint :  std_logic_vector(40 downto 0);
signal M :  std_logic_vector(40 downto 0);
signal Rtmp :  std_logic_vector(40 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(40 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_17x24_F50_uid28
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x24_F50_uid28 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(40 downto 0)   );
end entity;

architecture arch of DSPBlock_17x24_F50_uid28 is
signal Mint :  std_logic_vector(40 downto 0);
signal M :  std_logic_vector(40 downto 0);
signal Rtmp :  std_logic_vector(40 downto 0);
begin
   Mint <= std_logic_vector(unsigned(X) * unsigned(Y)); -- multiplier
   M <= Mint(40 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_10x24_F50_uid30
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_10x24_F50_uid30 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : in  std_logic_vector(23 downto 0);
          R : out  std_logic_vector(33 downto 0)   );
end entity;

architecture arch of DSPBlock_10x24_F50_uid30 is
signal Mint :  std_logic_vector(34 downto 0);
signal M :  std_logic_vector(33 downto 0);
signal Rtmp :  std_logic_vector(33 downto 0);
begin
   Mint <= std_logic_vector(signed(X) * signed('0' & Y)); -- multiplier
   M <= Mint(33 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_17x13_F50_uid32
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x13_F50_uid32 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(12 downto 0);
          R : out  std_logic_vector(29 downto 0)   );
end entity;

architecture arch of DSPBlock_17x13_F50_uid32 is
signal Mint :  std_logic_vector(30 downto 0);
signal M :  std_logic_vector(29 downto 0);
signal Rtmp :  std_logic_vector(29 downto 0);
begin
   Mint <= std_logic_vector(signed('0' & X) * signed(Y)); -- multiplier
   M <= Mint(29 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_17x13_F50_uid34
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x13_F50_uid34 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(12 downto 0);
          R : out  std_logic_vector(29 downto 0)   );
end entity;

architecture arch of DSPBlock_17x13_F50_uid34 is
signal Mint :  std_logic_vector(30 downto 0);
signal M :  std_logic_vector(29 downto 0);
signal Rtmp :  std_logic_vector(29 downto 0);
begin
   Mint <= std_logic_vector(signed('0' & X) * signed(Y)); -- multiplier
   M <= Mint(29 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_17x13_F50_uid36
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_17x13_F50_uid36 is
    port (clk : in std_logic;
          X : in  std_logic_vector(16 downto 0);
          Y : in  std_logic_vector(12 downto 0);
          R : out  std_logic_vector(29 downto 0)   );
end entity;

architecture arch of DSPBlock_17x13_F50_uid36 is
signal Mint :  std_logic_vector(30 downto 0);
signal M :  std_logic_vector(29 downto 0);
signal Rtmp :  std_logic_vector(29 downto 0);
begin
   Mint <= std_logic_vector(signed('0' & X) * signed(Y)); -- multiplier
   M <= Mint(29 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          DSPBlock_10x13_F50_uid38
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: 
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity DSPBlock_10x13_F50_uid38 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : in  std_logic_vector(12 downto 0);
          R : out  std_logic_vector(22 downto 0)   );
end entity;

architecture arch of DSPBlock_10x13_F50_uid38 is
signal Mint :  std_logic_vector(22 downto 0);
signal M :  std_logic_vector(22 downto 0);
signal Rtmp :  std_logic_vector(22 downto 0);
begin
   Mint <= std_logic_vector(signed(X) * signed(Y)); -- multiplier
   M <= Mint(22 downto 0);
   Rtmp <= M;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_100_F50_uid443
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_100_F50_uid443 is
    port (clk : in std_logic;
          X : in  std_logic_vector(99 downto 0);
          Y : in  std_logic_vector(99 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(99 downto 0)   );
end entity;

architecture arch of IntAdder_100_F50_uid443 is
signal Rtmp :  std_logic_vector(99 downto 0);
begin
   Rtmp <= X + Y + Cin;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                          IntMultiplier_F50_uid122
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Martin Kumm, Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_F50_uid122 is
    port (clk : in std_logic;
          X : in  std_logic_vector(60 downto 0);
          Y : in  std_logic_vector(60 downto 0);
          R : out  std_logic_vector(121 downto 0)   );
end entity;

architecture arch of IntMultiplier_F50_uid122 is
   component DSPBlock_17x24_F50_uid16 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_F50_uid18 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_F50_uid20 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_10x24_F50_uid22 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(33 downto 0)   );
   end component;

   component DSPBlock_17x24_F50_uid24 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_F50_uid26 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_17x24_F50_uid28 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(40 downto 0)   );
   end component;

   component DSPBlock_10x24_F50_uid30 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(33 downto 0)   );
   end component;

   component DSPBlock_17x13_F50_uid32 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(12 downto 0);
             R : out  std_logic_vector(29 downto 0)   );
   end component;

   component DSPBlock_17x13_F50_uid34 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(12 downto 0);
             R : out  std_logic_vector(29 downto 0)   );
   end component;

   component DSPBlock_17x13_F50_uid36 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(16 downto 0);
             Y : in  std_logic_vector(12 downto 0);
             R : out  std_logic_vector(29 downto 0)   );
   end component;

   component DSPBlock_10x13_F50_uid38 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : in  std_logic_vector(12 downto 0);
             R : out  std_logic_vector(22 downto 0)   );
   end component;

   component Compressor_23_3_F50_uid41 is
      port ( X1 : in  std_logic_vector(1 downto 0);
             X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2_F50_uid49 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

   component Compressor_14_3_F50_uid63 is
      port ( X1 : in  std_logic_vector(0 downto 0);
             X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_6_3_F50_uid99 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component IntAdder_100_F50_uid443 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(99 downto 0);
             Y : in  std_logic_vector(99 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(99 downto 0)   );
   end component;

signal XX_m13 :  std_logic_vector(60 downto 0);
signal YY_m13 :  std_logic_vector(60 downto 0);
signal tile_0_X :  std_logic_vector(16 downto 0);
signal tile_0_Y :  std_logic_vector(23 downto 0);
signal tile_0_output :  std_logic_vector(40 downto 0);
signal tile_0_filtered_output :  unsigned(40-0 downto 0);
signal bh14_w0_0 :  std_logic;
signal bh14_w1_0 :  std_logic;
signal bh14_w2_0 :  std_logic;
signal bh14_w3_0 :  std_logic;
signal bh14_w4_0 :  std_logic;
signal bh14_w5_0 :  std_logic;
signal bh14_w6_0 :  std_logic;
signal bh14_w7_0 :  std_logic;
signal bh14_w8_0 :  std_logic;
signal bh14_w9_0 :  std_logic;
signal bh14_w10_0 :  std_logic;
signal bh14_w11_0 :  std_logic;
signal bh14_w12_0 :  std_logic;
signal bh14_w13_0 :  std_logic;
signal bh14_w14_0 :  std_logic;
signal bh14_w15_0 :  std_logic;
signal bh14_w16_0 :  std_logic;
signal bh14_w17_0 :  std_logic;
signal bh14_w18_0 :  std_logic;
signal bh14_w19_0 :  std_logic;
signal bh14_w20_0 :  std_logic;
signal bh14_w21_0 :  std_logic;
signal bh14_w22_0 :  std_logic;
signal bh14_w23_0 :  std_logic;
signal bh14_w24_0 :  std_logic;
signal bh14_w25_0 :  std_logic;
signal bh14_w26_0 :  std_logic;
signal bh14_w27_0 :  std_logic;
signal bh14_w28_0 :  std_logic;
signal bh14_w29_0 :  std_logic;
signal bh14_w30_0 :  std_logic;
signal bh14_w31_0 :  std_logic;
signal bh14_w32_0 :  std_logic;
signal bh14_w33_0 :  std_logic;
signal bh14_w34_0 :  std_logic;
signal bh14_w35_0 :  std_logic;
signal bh14_w36_0 :  std_logic;
signal bh14_w37_0 :  std_logic;
signal bh14_w38_0 :  std_logic;
signal bh14_w39_0 :  std_logic;
signal bh14_w40_0 :  std_logic;
signal tile_1_X :  std_logic_vector(16 downto 0);
signal tile_1_Y :  std_logic_vector(23 downto 0);
signal tile_1_output :  std_logic_vector(40 downto 0);
signal tile_1_filtered_output :  unsigned(40-0 downto 0);
signal bh14_w17_1 :  std_logic;
signal bh14_w18_1 :  std_logic;
signal bh14_w19_1 :  std_logic;
signal bh14_w20_1 :  std_logic;
signal bh14_w21_1 :  std_logic;
signal bh14_w22_1 :  std_logic;
signal bh14_w23_1 :  std_logic;
signal bh14_w24_1 :  std_logic;
signal bh14_w25_1 :  std_logic;
signal bh14_w26_1 :  std_logic;
signal bh14_w27_1 :  std_logic;
signal bh14_w28_1 :  std_logic;
signal bh14_w29_1 :  std_logic;
signal bh14_w30_1 :  std_logic;
signal bh14_w31_1 :  std_logic;
signal bh14_w32_1 :  std_logic;
signal bh14_w33_1 :  std_logic;
signal bh14_w34_1 :  std_logic;
signal bh14_w35_1 :  std_logic;
signal bh14_w36_1 :  std_logic;
signal bh14_w37_1 :  std_logic;
signal bh14_w38_1 :  std_logic;
signal bh14_w39_1 :  std_logic;
signal bh14_w40_1 :  std_logic;
signal bh14_w41_0 :  std_logic;
signal bh14_w42_0 :  std_logic;
signal bh14_w43_0 :  std_logic;
signal bh14_w44_0 :  std_logic;
signal bh14_w45_0 :  std_logic;
signal bh14_w46_0 :  std_logic;
signal bh14_w47_0 :  std_logic;
signal bh14_w48_0 :  std_logic;
signal bh14_w49_0 :  std_logic;
signal bh14_w50_0 :  std_logic;
signal bh14_w51_0 :  std_logic;
signal bh14_w52_0 :  std_logic;
signal bh14_w53_0 :  std_logic;
signal bh14_w54_0 :  std_logic;
signal bh14_w55_0 :  std_logic;
signal bh14_w56_0 :  std_logic;
signal bh14_w57_0 :  std_logic;
signal tile_2_X :  std_logic_vector(16 downto 0);
signal tile_2_Y :  std_logic_vector(23 downto 0);
signal tile_2_output :  std_logic_vector(40 downto 0);
signal tile_2_filtered_output :  unsigned(40-0 downto 0);
signal bh14_w34_2 :  std_logic;
signal bh14_w35_2 :  std_logic;
signal bh14_w36_2 :  std_logic;
signal bh14_w37_2 :  std_logic;
signal bh14_w38_2 :  std_logic;
signal bh14_w39_2 :  std_logic;
signal bh14_w40_2 :  std_logic;
signal bh14_w41_1 :  std_logic;
signal bh14_w42_1 :  std_logic;
signal bh14_w43_1 :  std_logic;
signal bh14_w44_1 :  std_logic;
signal bh14_w45_1 :  std_logic;
signal bh14_w46_1 :  std_logic;
signal bh14_w47_1 :  std_logic;
signal bh14_w48_1 :  std_logic;
signal bh14_w49_1 :  std_logic;
signal bh14_w50_1 :  std_logic;
signal bh14_w51_1 :  std_logic;
signal bh14_w52_1 :  std_logic;
signal bh14_w53_1 :  std_logic;
signal bh14_w54_1 :  std_logic;
signal bh14_w55_1 :  std_logic;
signal bh14_w56_1 :  std_logic;
signal bh14_w57_1 :  std_logic;
signal bh14_w58_0 :  std_logic;
signal bh14_w59_0 :  std_logic;
signal bh14_w60_0 :  std_logic;
signal bh14_w61_0 :  std_logic;
signal bh14_w62_0 :  std_logic;
signal bh14_w63_0 :  std_logic;
signal bh14_w64_0 :  std_logic;
signal bh14_w65_0 :  std_logic;
signal bh14_w66_0 :  std_logic;
signal bh14_w67_0 :  std_logic;
signal bh14_w68_0 :  std_logic;
signal bh14_w69_0 :  std_logic;
signal bh14_w70_0 :  std_logic;
signal bh14_w71_0 :  std_logic;
signal bh14_w72_0 :  std_logic;
signal bh14_w73_0 :  std_logic;
signal bh14_w74_0 :  std_logic;
signal tile_3_X :  std_logic_vector(9 downto 0);
signal tile_3_Y :  std_logic_vector(23 downto 0);
signal tile_3_output :  std_logic_vector(33 downto 0);
signal tile_3_filtered_output :  signed(33-0 downto 0);
signal bh14_w51_2 :  std_logic;
signal bh14_w52_2 :  std_logic;
signal bh14_w53_2 :  std_logic;
signal bh14_w54_2 :  std_logic;
signal bh14_w55_2 :  std_logic;
signal bh14_w56_2 :  std_logic;
signal bh14_w57_2 :  std_logic;
signal bh14_w58_1 :  std_logic;
signal bh14_w59_1 :  std_logic;
signal bh14_w60_1 :  std_logic;
signal bh14_w61_1 :  std_logic;
signal bh14_w62_1 :  std_logic;
signal bh14_w63_1 :  std_logic;
signal bh14_w64_1 :  std_logic;
signal bh14_w65_1 :  std_logic;
signal bh14_w66_1 :  std_logic;
signal bh14_w67_1 :  std_logic;
signal bh14_w68_1 :  std_logic;
signal bh14_w69_1 :  std_logic;
signal bh14_w70_1 :  std_logic;
signal bh14_w71_1 :  std_logic;
signal bh14_w72_1 :  std_logic;
signal bh14_w73_1 :  std_logic;
signal bh14_w74_1 :  std_logic;
signal bh14_w75_0 :  std_logic;
signal bh14_w76_0 :  std_logic;
signal bh14_w77_0 :  std_logic;
signal bh14_w78_0 :  std_logic;
signal bh14_w79_0 :  std_logic;
signal bh14_w80_0 :  std_logic;
signal bh14_w81_0 :  std_logic;
signal bh14_w82_0 :  std_logic;
signal bh14_w83_0 :  std_logic;
signal bh14_w84_0 :  std_logic;
signal tile_4_X :  std_logic_vector(16 downto 0);
signal tile_4_Y :  std_logic_vector(23 downto 0);
signal tile_4_output :  std_logic_vector(40 downto 0);
signal tile_4_filtered_output :  unsigned(40-0 downto 0);
signal bh14_w24_2 :  std_logic;
signal bh14_w25_2 :  std_logic;
signal bh14_w26_2 :  std_logic;
signal bh14_w27_2 :  std_logic;
signal bh14_w28_2 :  std_logic;
signal bh14_w29_2 :  std_logic;
signal bh14_w30_2 :  std_logic;
signal bh14_w31_2 :  std_logic;
signal bh14_w32_2 :  std_logic;
signal bh14_w33_2 :  std_logic;
signal bh14_w34_3 :  std_logic;
signal bh14_w35_3 :  std_logic;
signal bh14_w36_3 :  std_logic;
signal bh14_w37_3 :  std_logic;
signal bh14_w38_3 :  std_logic;
signal bh14_w39_3 :  std_logic;
signal bh14_w40_3 :  std_logic;
signal bh14_w41_2 :  std_logic;
signal bh14_w42_2 :  std_logic;
signal bh14_w43_2 :  std_logic;
signal bh14_w44_2 :  std_logic;
signal bh14_w45_2 :  std_logic;
signal bh14_w46_2 :  std_logic;
signal bh14_w47_2 :  std_logic;
signal bh14_w48_2 :  std_logic;
signal bh14_w49_2 :  std_logic;
signal bh14_w50_2 :  std_logic;
signal bh14_w51_3 :  std_logic;
signal bh14_w52_3 :  std_logic;
signal bh14_w53_3 :  std_logic;
signal bh14_w54_3 :  std_logic;
signal bh14_w55_3 :  std_logic;
signal bh14_w56_3 :  std_logic;
signal bh14_w57_3 :  std_logic;
signal bh14_w58_2 :  std_logic;
signal bh14_w59_2 :  std_logic;
signal bh14_w60_2 :  std_logic;
signal bh14_w61_2 :  std_logic;
signal bh14_w62_2 :  std_logic;
signal bh14_w63_2 :  std_logic;
signal bh14_w64_2 :  std_logic;
signal tile_5_X :  std_logic_vector(16 downto 0);
signal tile_5_Y :  std_logic_vector(23 downto 0);
signal tile_5_output :  std_logic_vector(40 downto 0);
signal tile_5_filtered_output :  unsigned(40-0 downto 0);
signal bh14_w41_3 :  std_logic;
signal bh14_w42_3 :  std_logic;
signal bh14_w43_3 :  std_logic;
signal bh14_w44_3 :  std_logic;
signal bh14_w45_3 :  std_logic;
signal bh14_w46_3 :  std_logic;
signal bh14_w47_3 :  std_logic;
signal bh14_w48_3 :  std_logic;
signal bh14_w49_3 :  std_logic;
signal bh14_w50_3 :  std_logic;
signal bh14_w51_4 :  std_logic;
signal bh14_w52_4 :  std_logic;
signal bh14_w53_4 :  std_logic;
signal bh14_w54_4 :  std_logic;
signal bh14_w55_4 :  std_logic;
signal bh14_w56_4 :  std_logic;
signal bh14_w57_4 :  std_logic;
signal bh14_w58_3 :  std_logic;
signal bh14_w59_3 :  std_logic;
signal bh14_w60_3 :  std_logic;
signal bh14_w61_3 :  std_logic;
signal bh14_w62_3 :  std_logic;
signal bh14_w63_3 :  std_logic;
signal bh14_w64_3 :  std_logic;
signal bh14_w65_2 :  std_logic;
signal bh14_w66_2 :  std_logic;
signal bh14_w67_2 :  std_logic;
signal bh14_w68_2 :  std_logic;
signal bh14_w69_2 :  std_logic;
signal bh14_w70_2 :  std_logic;
signal bh14_w71_2 :  std_logic;
signal bh14_w72_2 :  std_logic;
signal bh14_w73_2 :  std_logic;
signal bh14_w74_2 :  std_logic;
signal bh14_w75_1 :  std_logic;
signal bh14_w76_1 :  std_logic;
signal bh14_w77_1 :  std_logic;
signal bh14_w78_1 :  std_logic;
signal bh14_w79_1 :  std_logic;
signal bh14_w80_1 :  std_logic;
signal bh14_w81_1 :  std_logic;
signal tile_6_X :  std_logic_vector(16 downto 0);
signal tile_6_Y :  std_logic_vector(23 downto 0);
signal tile_6_output :  std_logic_vector(40 downto 0);
signal tile_6_filtered_output :  unsigned(40-0 downto 0);
signal bh14_w58_4 :  std_logic;
signal bh14_w59_4 :  std_logic;
signal bh14_w60_4 :  std_logic;
signal bh14_w61_4 :  std_logic;
signal bh14_w62_4 :  std_logic;
signal bh14_w63_4 :  std_logic;
signal bh14_w64_4 :  std_logic;
signal bh14_w65_3 :  std_logic;
signal bh14_w66_3 :  std_logic;
signal bh14_w67_3 :  std_logic;
signal bh14_w68_3 :  std_logic;
signal bh14_w69_3 :  std_logic;
signal bh14_w70_3 :  std_logic;
signal bh14_w71_3 :  std_logic;
signal bh14_w72_3 :  std_logic;
signal bh14_w73_3 :  std_logic;
signal bh14_w74_3 :  std_logic;
signal bh14_w75_2 :  std_logic;
signal bh14_w76_2 :  std_logic;
signal bh14_w77_2 :  std_logic;
signal bh14_w78_2 :  std_logic;
signal bh14_w79_2 :  std_logic;
signal bh14_w80_2 :  std_logic;
signal bh14_w81_2 :  std_logic;
signal bh14_w82_1 :  std_logic;
signal bh14_w83_1 :  std_logic;
signal bh14_w84_1 :  std_logic;
signal bh14_w85_0 :  std_logic;
signal bh14_w86_0 :  std_logic;
signal bh14_w87_0 :  std_logic;
signal bh14_w88_0 :  std_logic;
signal bh14_w89_0 :  std_logic;
signal bh14_w90_0 :  std_logic;
signal bh14_w91_0 :  std_logic;
signal bh14_w92_0 :  std_logic;
signal bh14_w93_0 :  std_logic;
signal bh14_w94_0 :  std_logic;
signal bh14_w95_0 :  std_logic;
signal bh14_w96_0 :  std_logic;
signal bh14_w97_0 :  std_logic;
signal bh14_w98_0 :  std_logic;
signal tile_7_X :  std_logic_vector(9 downto 0);
signal tile_7_Y :  std_logic_vector(23 downto 0);
signal tile_7_output :  std_logic_vector(33 downto 0);
signal tile_7_filtered_output :  signed(33-0 downto 0);
signal bh14_w75_3 :  std_logic;
signal bh14_w76_3 :  std_logic;
signal bh14_w77_3 :  std_logic;
signal bh14_w78_3 :  std_logic;
signal bh14_w79_3 :  std_logic;
signal bh14_w80_3 :  std_logic;
signal bh14_w81_3 :  std_logic;
signal bh14_w82_2 :  std_logic;
signal bh14_w83_2 :  std_logic;
signal bh14_w84_2 :  std_logic;
signal bh14_w85_1 :  std_logic;
signal bh14_w86_1 :  std_logic;
signal bh14_w87_1 :  std_logic;
signal bh14_w88_1 :  std_logic;
signal bh14_w89_1 :  std_logic;
signal bh14_w90_1 :  std_logic;
signal bh14_w91_1 :  std_logic;
signal bh14_w92_1 :  std_logic;
signal bh14_w93_1 :  std_logic;
signal bh14_w94_1 :  std_logic;
signal bh14_w95_1 :  std_logic;
signal bh14_w96_1 :  std_logic;
signal bh14_w97_1 :  std_logic;
signal bh14_w98_1 :  std_logic;
signal bh14_w99_0 :  std_logic;
signal bh14_w100_0 :  std_logic;
signal bh14_w101_0 :  std_logic;
signal bh14_w102_0 :  std_logic;
signal bh14_w103_0 :  std_logic;
signal bh14_w104_0 :  std_logic;
signal bh14_w105_0 :  std_logic;
signal bh14_w106_0 :  std_logic;
signal bh14_w107_0 :  std_logic;
signal bh14_w108_0 :  std_logic;
signal tile_8_X :  std_logic_vector(16 downto 0);
signal tile_8_Y :  std_logic_vector(12 downto 0);
signal tile_8_output :  std_logic_vector(29 downto 0);
signal tile_8_filtered_output :  signed(29-0 downto 0);
signal bh14_w48_4 :  std_logic;
signal bh14_w49_4 :  std_logic;
signal bh14_w50_4 :  std_logic;
signal bh14_w51_5 :  std_logic;
signal bh14_w52_5 :  std_logic;
signal bh14_w53_5 :  std_logic;
signal bh14_w54_5 :  std_logic;
signal bh14_w55_5 :  std_logic;
signal bh14_w56_5 :  std_logic;
signal bh14_w57_5 :  std_logic;
signal bh14_w58_5 :  std_logic;
signal bh14_w59_5 :  std_logic;
signal bh14_w60_5 :  std_logic;
signal bh14_w61_5 :  std_logic;
signal bh14_w62_5 :  std_logic;
signal bh14_w63_5 :  std_logic;
signal bh14_w64_5 :  std_logic;
signal bh14_w65_4 :  std_logic;
signal bh14_w66_4 :  std_logic;
signal bh14_w67_4 :  std_logic;
signal bh14_w68_4 :  std_logic;
signal bh14_w69_4 :  std_logic;
signal bh14_w70_4 :  std_logic;
signal bh14_w71_4 :  std_logic;
signal bh14_w72_4 :  std_logic;
signal bh14_w73_4 :  std_logic;
signal bh14_w74_4 :  std_logic;
signal bh14_w75_4 :  std_logic;
signal bh14_w76_4 :  std_logic;
signal bh14_w77_4 :  std_logic;
signal tile_9_X :  std_logic_vector(16 downto 0);
signal tile_9_Y :  std_logic_vector(12 downto 0);
signal tile_9_output :  std_logic_vector(29 downto 0);
signal tile_9_filtered_output :  signed(29-0 downto 0);
signal bh14_w65_5 :  std_logic;
signal bh14_w66_5 :  std_logic;
signal bh14_w67_5 :  std_logic;
signal bh14_w68_5 :  std_logic;
signal bh14_w69_5 :  std_logic;
signal bh14_w70_5 :  std_logic;
signal bh14_w71_5 :  std_logic;
signal bh14_w72_5 :  std_logic;
signal bh14_w73_5 :  std_logic;
signal bh14_w74_5 :  std_logic;
signal bh14_w75_5 :  std_logic;
signal bh14_w76_5 :  std_logic;
signal bh14_w77_5 :  std_logic;
signal bh14_w78_4 :  std_logic;
signal bh14_w79_4 :  std_logic;
signal bh14_w80_4 :  std_logic;
signal bh14_w81_4 :  std_logic;
signal bh14_w82_3 :  std_logic;
signal bh14_w83_3 :  std_logic;
signal bh14_w84_3 :  std_logic;
signal bh14_w85_2 :  std_logic;
signal bh14_w86_2 :  std_logic;
signal bh14_w87_2 :  std_logic;
signal bh14_w88_2 :  std_logic;
signal bh14_w89_2 :  std_logic;
signal bh14_w90_2 :  std_logic;
signal bh14_w91_2 :  std_logic;
signal bh14_w92_2 :  std_logic;
signal bh14_w93_2 :  std_logic;
signal bh14_w94_2 :  std_logic;
signal tile_10_X :  std_logic_vector(16 downto 0);
signal tile_10_Y :  std_logic_vector(12 downto 0);
signal tile_10_output :  std_logic_vector(29 downto 0);
signal tile_10_filtered_output :  signed(29-0 downto 0);
signal bh14_w82_4 :  std_logic;
signal bh14_w83_4 :  std_logic;
signal bh14_w84_4 :  std_logic;
signal bh14_w85_3 :  std_logic;
signal bh14_w86_3 :  std_logic;
signal bh14_w87_3 :  std_logic;
signal bh14_w88_3 :  std_logic;
signal bh14_w89_3 :  std_logic;
signal bh14_w90_3 :  std_logic;
signal bh14_w91_3 :  std_logic;
signal bh14_w92_3 :  std_logic;
signal bh14_w93_3 :  std_logic;
signal bh14_w94_3 :  std_logic;
signal bh14_w95_2 :  std_logic;
signal bh14_w96_2 :  std_logic;
signal bh14_w97_2 :  std_logic;
signal bh14_w98_2 :  std_logic;
signal bh14_w99_1 :  std_logic;
signal bh14_w100_1 :  std_logic;
signal bh14_w101_1 :  std_logic;
signal bh14_w102_1 :  std_logic;
signal bh14_w103_1 :  std_logic;
signal bh14_w104_1 :  std_logic;
signal bh14_w105_1 :  std_logic;
signal bh14_w106_1 :  std_logic;
signal bh14_w107_1 :  std_logic;
signal bh14_w108_1 :  std_logic;
signal bh14_w109_0 :  std_logic;
signal bh14_w110_0 :  std_logic;
signal bh14_w111_0 :  std_logic;
signal tile_11_X :  std_logic_vector(9 downto 0);
signal tile_11_Y :  std_logic_vector(12 downto 0);
signal tile_11_output :  std_logic_vector(22 downto 0);
signal tile_11_filtered_output :  signed(22-0 downto 0);
signal bh14_w99_2 :  std_logic;
signal bh14_w100_2 :  std_logic;
signal bh14_w101_2 :  std_logic;
signal bh14_w102_2 :  std_logic;
signal bh14_w103_2 :  std_logic;
signal bh14_w104_2 :  std_logic;
signal bh14_w105_2 :  std_logic;
signal bh14_w106_2 :  std_logic;
signal bh14_w107_2 :  std_logic;
signal bh14_w108_2 :  std_logic;
signal bh14_w109_1 :  std_logic;
signal bh14_w110_1 :  std_logic;
signal bh14_w111_1 :  std_logic;
signal bh14_w112_0 :  std_logic;
signal bh14_w113_0 :  std_logic;
signal bh14_w114_0 :  std_logic;
signal bh14_w115_0 :  std_logic;
signal bh14_w116_0 :  std_logic;
signal bh14_w117_0 :  std_logic;
signal bh14_w118_0 :  std_logic;
signal bh14_w119_0 :  std_logic;
signal bh14_w120_0 :  std_logic;
signal bh14_w121_0 :  std_logic;
signal bh14_w77_6 :  std_logic;
signal bh14_w78_5 :  std_logic;
signal bh14_w79_5 :  std_logic;
signal bh14_w80_5 :  std_logic;
signal bh14_w81_5 :  std_logic;
signal bh14_w82_5 :  std_logic;
signal bh14_w83_5 :  std_logic;
signal bh14_w85_4 :  std_logic;
signal bh14_w86_4 :  std_logic;
signal bh14_w87_4 :  std_logic;
signal bh14_w88_4 :  std_logic;
signal bh14_w89_4 :  std_logic;
signal bh14_w90_4 :  std_logic;
signal bh14_w91_4 :  std_logic;
signal bh14_w92_4 :  std_logic;
signal bh14_w93_4 :  std_logic;
signal bh14_w95_3 :  std_logic;
signal bh14_w96_3 :  std_logic;
signal bh14_w97_3 :  std_logic;
signal bh14_w98_3 :  std_logic;
signal bh14_w99_3 :  std_logic;
signal bh14_w100_3 :  std_logic;
signal bh14_w101_3 :  std_logic;
signal bh14_w102_3 :  std_logic;
signal bh14_w103_3 :  std_logic;
signal bh14_w104_3 :  std_logic;
signal bh14_w105_3 :  std_logic;
signal bh14_w106_3 :  std_logic;
signal bh14_w107_3 :  std_logic;
signal bh14_w109_2 :  std_logic;
signal bh14_w110_2 :  std_logic;
signal bh14_w112_1 :  std_logic;
signal bh14_w113_1 :  std_logic;
signal bh14_w114_1 :  std_logic;
signal bh14_w115_1 :  std_logic;
signal bh14_w116_1 :  std_logic;
signal bh14_w117_1 :  std_logic;
signal bh14_w118_1 :  std_logic;
signal bh14_w119_1 :  std_logic;
signal bh14_w120_1 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid42_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid42_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid42_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid42_Out0_copy43 :  std_logic_vector(2 downto 0);
signal bh14_w17_2 :  std_logic;
signal bh14_w18_2 :  std_logic;
signal bh14_w19_2 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid44_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid44_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid44_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid44_Out0_copy45 :  std_logic_vector(2 downto 0);
signal bh14_w19_3 :  std_logic;
signal bh14_w20_2 :  std_logic;
signal bh14_w21_2 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid46_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid46_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid46_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid46_Out0_copy47 :  std_logic_vector(2 downto 0);
signal bh14_w21_3 :  std_logic;
signal bh14_w22_2 :  std_logic;
signal bh14_w23_2 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid50_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid50_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid50_Out0_copy51 :  std_logic_vector(1 downto 0);
signal bh14_w23_3 :  std_logic;
signal bh14_w24_3 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid52_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid52_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid52_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid52_Out0_copy53 :  std_logic_vector(2 downto 0);
signal bh14_w24_4 :  std_logic;
signal bh14_w25_3 :  std_logic;
signal bh14_w26_3 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid54_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid54_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid54_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid54_Out0_copy55 :  std_logic_vector(2 downto 0);
signal bh14_w26_4 :  std_logic;
signal bh14_w27_3 :  std_logic;
signal bh14_w28_3 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid56_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid56_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid56_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid56_Out0_copy57 :  std_logic_vector(2 downto 0);
signal bh14_w28_4 :  std_logic;
signal bh14_w29_3 :  std_logic;
signal bh14_w30_3 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid58_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid58_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid58_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid58_Out0_copy59 :  std_logic_vector(2 downto 0);
signal bh14_w30_4 :  std_logic;
signal bh14_w31_3 :  std_logic;
signal bh14_w32_3 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid60_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid60_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid60_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid60_Out0_copy61 :  std_logic_vector(2 downto 0);
signal bh14_w32_4 :  std_logic;
signal bh14_w33_3 :  std_logic;
signal bh14_w34_4 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid64_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid64_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid64_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid64_Out0_copy65 :  std_logic_vector(2 downto 0);
signal bh14_w34_5 :  std_logic;
signal bh14_w35_4 :  std_logic;
signal bh14_w36_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid66_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid66_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid66_Out0_copy67 :  std_logic_vector(1 downto 0);
signal bh14_w35_5 :  std_logic;
signal bh14_w36_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid68_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid68_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid68_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid68_Out0_copy69 :  std_logic_vector(2 downto 0);
signal bh14_w36_6 :  std_logic;
signal bh14_w37_4 :  std_logic;
signal bh14_w38_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid70_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid70_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid70_Out0_copy71 :  std_logic_vector(1 downto 0);
signal bh14_w37_5 :  std_logic;
signal bh14_w38_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid72_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid72_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid72_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid72_Out0_copy73 :  std_logic_vector(2 downto 0);
signal bh14_w38_6 :  std_logic;
signal bh14_w39_4 :  std_logic;
signal bh14_w40_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid74_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid74_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid74_Out0_copy75 :  std_logic_vector(1 downto 0);
signal bh14_w39_5 :  std_logic;
signal bh14_w40_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid76_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid76_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid76_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid76_Out0_copy77 :  std_logic_vector(2 downto 0);
signal bh14_w40_6 :  std_logic;
signal bh14_w41_4 :  std_logic;
signal bh14_w42_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid78_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid78_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid78_Out0_copy79 :  std_logic_vector(1 downto 0);
signal bh14_w41_5 :  std_logic;
signal bh14_w42_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid80_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid80_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid80_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid80_Out0_copy81 :  std_logic_vector(2 downto 0);
signal bh14_w42_6 :  std_logic;
signal bh14_w43_4 :  std_logic;
signal bh14_w44_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid82_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid82_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid82_Out0_copy83 :  std_logic_vector(1 downto 0);
signal bh14_w43_5 :  std_logic;
signal bh14_w44_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid84_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid84_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid84_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid84_Out0_copy85 :  std_logic_vector(2 downto 0);
signal bh14_w44_6 :  std_logic;
signal bh14_w45_4 :  std_logic;
signal bh14_w46_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid86_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid86_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid86_Out0_copy87 :  std_logic_vector(1 downto 0);
signal bh14_w45_5 :  std_logic;
signal bh14_w46_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid88_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid88_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid88_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid88_Out0_copy89 :  std_logic_vector(2 downto 0);
signal bh14_w46_6 :  std_logic;
signal bh14_w47_4 :  std_logic;
signal bh14_w48_5 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid90_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid90_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid90_Out0_copy91 :  std_logic_vector(1 downto 0);
signal bh14_w47_5 :  std_logic;
signal bh14_w48_6 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid92_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid92_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid92_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid92_Out0_copy93 :  std_logic_vector(2 downto 0);
signal bh14_w48_7 :  std_logic;
signal bh14_w49_5 :  std_logic;
signal bh14_w50_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid94_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid94_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid94_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid94_Out0_copy95 :  std_logic_vector(2 downto 0);
signal bh14_w49_6 :  std_logic;
signal bh14_w50_6 :  std_logic;
signal bh14_w51_6 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid96_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid96_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid96_Out0_copy97 :  std_logic_vector(1 downto 0);
signal bh14_w50_7 :  std_logic;
signal bh14_w51_7 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid100_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid100_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid100_Out0_copy101 :  std_logic_vector(2 downto 0);
signal bh14_w51_8 :  std_logic;
signal bh14_w52_6 :  std_logic;
signal bh14_w53_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid102_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid102_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid102_Out0_copy103 :  std_logic_vector(2 downto 0);
signal bh14_w52_7 :  std_logic;
signal bh14_w53_7 :  std_logic;
signal bh14_w54_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid104_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid104_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid104_Out0_copy105 :  std_logic_vector(2 downto 0);
signal bh14_w53_8 :  std_logic;
signal bh14_w54_7 :  std_logic;
signal bh14_w55_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid106_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid106_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid106_Out0_copy107 :  std_logic_vector(2 downto 0);
signal bh14_w54_8 :  std_logic;
signal bh14_w55_7 :  std_logic;
signal bh14_w56_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid108_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid108_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid108_Out0_copy109 :  std_logic_vector(2 downto 0);
signal bh14_w55_8 :  std_logic;
signal bh14_w56_7 :  std_logic;
signal bh14_w57_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid110_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid110_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid110_Out0_copy111 :  std_logic_vector(2 downto 0);
signal bh14_w56_8 :  std_logic;
signal bh14_w57_7 :  std_logic;
signal bh14_w58_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid112_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid112_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid112_Out0_copy113 :  std_logic_vector(2 downto 0);
signal bh14_w57_8 :  std_logic;
signal bh14_w58_7 :  std_logic;
signal bh14_w59_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid114_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid114_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid114_Out0_copy115 :  std_logic_vector(2 downto 0);
signal bh14_w58_8 :  std_logic;
signal bh14_w59_7 :  std_logic;
signal bh14_w60_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid116_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid116_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid116_Out0_copy117 :  std_logic_vector(2 downto 0);
signal bh14_w59_8 :  std_logic;
signal bh14_w60_7 :  std_logic;
signal bh14_w61_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid118_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid118_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid118_Out0_copy119 :  std_logic_vector(2 downto 0);
signal bh14_w60_8 :  std_logic;
signal bh14_w61_7 :  std_logic;
signal bh14_w62_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid120_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid120_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid120_Out0_copy121 :  std_logic_vector(2 downto 0);
signal bh14_w61_8 :  std_logic;
signal bh14_w62_7 :  std_logic;
signal bh14_w63_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid122_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid122_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid122_Out0_copy123 :  std_logic_vector(2 downto 0);
signal bh14_w62_8 :  std_logic;
signal bh14_w63_7 :  std_logic;
signal bh14_w64_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid124_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid124_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid124_Out0_copy125 :  std_logic_vector(2 downto 0);
signal bh14_w63_8 :  std_logic;
signal bh14_w64_7 :  std_logic;
signal bh14_w65_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid126_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid126_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid126_Out0_copy127 :  std_logic_vector(2 downto 0);
signal bh14_w64_8 :  std_logic;
signal bh14_w65_7 :  std_logic;
signal bh14_w66_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid128_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid128_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid128_Out0_copy129 :  std_logic_vector(2 downto 0);
signal bh14_w65_8 :  std_logic;
signal bh14_w66_7 :  std_logic;
signal bh14_w67_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid130_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid130_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid130_Out0_copy131 :  std_logic_vector(2 downto 0);
signal bh14_w66_8 :  std_logic;
signal bh14_w67_7 :  std_logic;
signal bh14_w68_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid132_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid132_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid132_Out0_copy133 :  std_logic_vector(2 downto 0);
signal bh14_w67_8 :  std_logic;
signal bh14_w68_7 :  std_logic;
signal bh14_w69_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid134_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid134_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid134_Out0_copy135 :  std_logic_vector(2 downto 0);
signal bh14_w68_8 :  std_logic;
signal bh14_w69_7 :  std_logic;
signal bh14_w70_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid136_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid136_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid136_Out0_copy137 :  std_logic_vector(2 downto 0);
signal bh14_w69_8 :  std_logic;
signal bh14_w70_7 :  std_logic;
signal bh14_w71_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid138_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid138_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid138_Out0_copy139 :  std_logic_vector(2 downto 0);
signal bh14_w70_8 :  std_logic;
signal bh14_w71_7 :  std_logic;
signal bh14_w72_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid140_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid140_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid140_Out0_copy141 :  std_logic_vector(2 downto 0);
signal bh14_w71_8 :  std_logic;
signal bh14_w72_7 :  std_logic;
signal bh14_w73_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid142_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid142_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid142_Out0_copy143 :  std_logic_vector(2 downto 0);
signal bh14_w72_8 :  std_logic;
signal bh14_w73_7 :  std_logic;
signal bh14_w74_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid144_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid144_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid144_Out0_copy145 :  std_logic_vector(2 downto 0);
signal bh14_w73_8 :  std_logic;
signal bh14_w74_7 :  std_logic;
signal bh14_w75_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid146_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid146_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid146_Out0_copy147 :  std_logic_vector(2 downto 0);
signal bh14_w74_8 :  std_logic;
signal bh14_w75_7 :  std_logic;
signal bh14_w76_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid148_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid148_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid148_Out0_copy149 :  std_logic_vector(2 downto 0);
signal bh14_w75_8 :  std_logic;
signal bh14_w76_7 :  std_logic;
signal bh14_w77_7 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid150_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid150_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid150_Out0_copy151 :  std_logic_vector(2 downto 0);
signal bh14_w76_8 :  std_logic;
signal bh14_w77_8 :  std_logic;
signal bh14_w78_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid152_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid152_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid152_Out0_copy153 :  std_logic_vector(2 downto 0);
signal bh14_w77_9 :  std_logic;
signal bh14_w78_7 :  std_logic;
signal bh14_w79_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid154_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid154_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid154_Out0_copy155 :  std_logic_vector(2 downto 0);
signal bh14_w78_8 :  std_logic;
signal bh14_w79_7 :  std_logic;
signal bh14_w80_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid156_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid156_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid156_Out0_copy157 :  std_logic_vector(2 downto 0);
signal bh14_w79_8 :  std_logic;
signal bh14_w80_7 :  std_logic;
signal bh14_w81_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid158_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid158_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid158_Out0_copy159 :  std_logic_vector(2 downto 0);
signal bh14_w80_8 :  std_logic;
signal bh14_w81_7 :  std_logic;
signal bh14_w82_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid160_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid160_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid160_Out0_copy161 :  std_logic_vector(2 downto 0);
signal bh14_w81_8 :  std_logic;
signal bh14_w82_7 :  std_logic;
signal bh14_w83_6 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid162_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid162_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid162_Out0_copy163 :  std_logic_vector(2 downto 0);
signal bh14_w82_8 :  std_logic;
signal bh14_w83_7 :  std_logic;
signal bh14_w84_5 :  std_logic;
signal Compressor_6_3_F50_uid99_bh14_uid164_In0 :  std_logic_vector(5 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid164_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_6_3_F50_uid99_bh14_uid164_Out0_copy165 :  std_logic_vector(2 downto 0);
signal bh14_w83_8 :  std_logic;
signal bh14_w84_6 :  std_logic;
signal bh14_w85_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid166_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid166_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid166_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid166_Out0_copy167 :  std_logic_vector(2 downto 0);
signal bh14_w84_7 :  std_logic;
signal bh14_w85_6 :  std_logic;
signal bh14_w86_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid168_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid168_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid168_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid168_Out0_copy169 :  std_logic_vector(2 downto 0);
signal bh14_w85_7 :  std_logic;
signal bh14_w86_6 :  std_logic;
signal bh14_w87_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid170_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid170_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid170_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid170_Out0_copy171 :  std_logic_vector(2 downto 0);
signal bh14_w86_7 :  std_logic;
signal bh14_w87_6 :  std_logic;
signal bh14_w88_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid172_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid172_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid172_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid172_Out0_copy173 :  std_logic_vector(2 downto 0);
signal bh14_w87_7 :  std_logic;
signal bh14_w88_6 :  std_logic;
signal bh14_w89_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid174_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid174_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid174_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid174_Out0_copy175 :  std_logic_vector(2 downto 0);
signal bh14_w88_7 :  std_logic;
signal bh14_w89_6 :  std_logic;
signal bh14_w90_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid176_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid176_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid176_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid176_Out0_copy177 :  std_logic_vector(2 downto 0);
signal bh14_w89_7 :  std_logic;
signal bh14_w90_6 :  std_logic;
signal bh14_w91_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid178_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid178_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid178_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid178_Out0_copy179 :  std_logic_vector(2 downto 0);
signal bh14_w90_7 :  std_logic;
signal bh14_w91_6 :  std_logic;
signal bh14_w92_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid180_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid180_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid180_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid180_Out0_copy181 :  std_logic_vector(2 downto 0);
signal bh14_w91_7 :  std_logic;
signal bh14_w92_6 :  std_logic;
signal bh14_w93_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid182_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid182_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid182_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid182_Out0_copy183 :  std_logic_vector(2 downto 0);
signal bh14_w92_7 :  std_logic;
signal bh14_w93_6 :  std_logic;
signal bh14_w94_4 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid184_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid184_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid184_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid184_Out0_copy185 :  std_logic_vector(2 downto 0);
signal bh14_w93_7 :  std_logic;
signal bh14_w94_5 :  std_logic;
signal bh14_w95_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid186_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid186_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid186_Out0_copy187 :  std_logic_vector(1 downto 0);
signal bh14_w94_6 :  std_logic;
signal bh14_w95_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid188_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid188_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid188_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid188_Out0_copy189 :  std_logic_vector(2 downto 0);
signal bh14_w95_6 :  std_logic;
signal bh14_w96_4 :  std_logic;
signal bh14_w97_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid190_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid190_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid190_Out0_copy191 :  std_logic_vector(1 downto 0);
signal bh14_w96_5 :  std_logic;
signal bh14_w97_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid192_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid192_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid192_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid192_Out0_copy193 :  std_logic_vector(2 downto 0);
signal bh14_w97_6 :  std_logic;
signal bh14_w98_4 :  std_logic;
signal bh14_w99_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid194_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid194_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid194_Out0_copy195 :  std_logic_vector(1 downto 0);
signal bh14_w98_5 :  std_logic;
signal bh14_w99_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid196_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid196_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid196_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid196_Out0_copy197 :  std_logic_vector(2 downto 0);
signal bh14_w99_6 :  std_logic;
signal bh14_w100_4 :  std_logic;
signal bh14_w101_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid198_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid198_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid198_Out0_copy199 :  std_logic_vector(1 downto 0);
signal bh14_w100_5 :  std_logic;
signal bh14_w101_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid200_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid200_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid200_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid200_Out0_copy201 :  std_logic_vector(2 downto 0);
signal bh14_w101_6 :  std_logic;
signal bh14_w102_4 :  std_logic;
signal bh14_w103_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid202_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid202_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid202_Out0_copy203 :  std_logic_vector(1 downto 0);
signal bh14_w102_5 :  std_logic;
signal bh14_w103_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid204_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid204_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid204_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid204_Out0_copy205 :  std_logic_vector(2 downto 0);
signal bh14_w103_6 :  std_logic;
signal bh14_w104_4 :  std_logic;
signal bh14_w105_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid206_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid206_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid206_Out0_copy207 :  std_logic_vector(1 downto 0);
signal bh14_w104_5 :  std_logic;
signal bh14_w105_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid208_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid208_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid208_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid208_Out0_copy209 :  std_logic_vector(2 downto 0);
signal bh14_w105_6 :  std_logic;
signal bh14_w106_4 :  std_logic;
signal bh14_w107_4 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid210_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid210_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid210_Out0_copy211 :  std_logic_vector(1 downto 0);
signal bh14_w106_5 :  std_logic;
signal bh14_w107_5 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid212_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid212_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid212_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid212_Out0_copy213 :  std_logic_vector(2 downto 0);
signal bh14_w107_6 :  std_logic;
signal bh14_w108_3 :  std_logic;
signal bh14_w109_3 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid214_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid214_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid214_Out0_copy215 :  std_logic_vector(1 downto 0);
signal bh14_w108_4 :  std_logic;
signal bh14_w109_4 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid216_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid216_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid216_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid216_Out0_copy217 :  std_logic_vector(2 downto 0);
signal bh14_w109_5 :  std_logic;
signal bh14_w110_3 :  std_logic;
signal bh14_w111_2 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid218_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid218_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid218_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid218_Out0_copy219 :  std_logic_vector(2 downto 0);
signal bh14_w111_3 :  std_logic;
signal bh14_w112_2 :  std_logic;
signal bh14_w113_2 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid220_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid220_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid220_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid220_Out0_copy221 :  std_logic_vector(2 downto 0);
signal bh14_w113_3 :  std_logic;
signal bh14_w114_2 :  std_logic;
signal bh14_w115_2 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid222_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid222_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid222_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid222_Out0_copy223 :  std_logic_vector(2 downto 0);
signal bh14_w115_3 :  std_logic;
signal bh14_w116_2 :  std_logic;
signal bh14_w117_2 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid224_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid224_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid224_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid224_Out0_copy225 :  std_logic_vector(2 downto 0);
signal bh14_w117_3 :  std_logic;
signal bh14_w118_2 :  std_logic;
signal bh14_w119_2 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid226_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid226_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid226_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid226_Out0_copy227 :  std_logic_vector(2 downto 0);
signal bh14_w119_3 :  std_logic;
signal bh14_w120_2 :  std_logic;
signal bh14_w121_1 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid228_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid228_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid228_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid228_Out0_copy229 :  std_logic_vector(2 downto 0);
signal bh14_w19_4 :  std_logic;
signal bh14_w20_3 :  std_logic;
signal bh14_w21_4 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid230_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid230_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid230_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid230_Out0_copy231 :  std_logic_vector(2 downto 0);
signal bh14_w21_5 :  std_logic;
signal bh14_w22_3 :  std_logic;
signal bh14_w23_4 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid232_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid232_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid232_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid232_Out0_copy233 :  std_logic_vector(2 downto 0);
signal bh14_w23_5 :  std_logic;
signal bh14_w24_5 :  std_logic;
signal bh14_w25_4 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid234_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid234_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid234_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid234_Out0_copy235 :  std_logic_vector(2 downto 0);
signal bh14_w25_5 :  std_logic;
signal bh14_w26_5 :  std_logic;
signal bh14_w27_4 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid236_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid236_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid236_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid236_Out0_copy237 :  std_logic_vector(2 downto 0);
signal bh14_w27_5 :  std_logic;
signal bh14_w28_5 :  std_logic;
signal bh14_w29_4 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid238_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid238_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid238_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid238_Out0_copy239 :  std_logic_vector(2 downto 0);
signal bh14_w29_5 :  std_logic;
signal bh14_w30_5 :  std_logic;
signal bh14_w31_4 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid240_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid240_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid240_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid240_Out0_copy241 :  std_logic_vector(2 downto 0);
signal bh14_w31_5 :  std_logic;
signal bh14_w32_5 :  std_logic;
signal bh14_w33_4 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid242_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid242_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid242_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid242_Out0_copy243 :  std_logic_vector(2 downto 0);
signal bh14_w33_5 :  std_logic;
signal bh14_w34_6 :  std_logic;
signal bh14_w35_6 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid244_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid244_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid244_Out0_copy245 :  std_logic_vector(1 downto 0);
signal bh14_w35_7 :  std_logic;
signal bh14_w36_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid246_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid246_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid246_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid246_Out0_copy247 :  std_logic_vector(2 downto 0);
signal bh14_w36_8 :  std_logic;
signal bh14_w37_6 :  std_logic;
signal bh14_w38_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid248_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid248_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid248_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid248_Out0_copy249 :  std_logic_vector(2 downto 0);
signal bh14_w38_8 :  std_logic;
signal bh14_w39_6 :  std_logic;
signal bh14_w40_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid250_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid250_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid250_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid250_Out0_copy251 :  std_logic_vector(2 downto 0);
signal bh14_w40_8 :  std_logic;
signal bh14_w41_6 :  std_logic;
signal bh14_w42_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid252_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid252_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid252_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid252_Out0_copy253 :  std_logic_vector(2 downto 0);
signal bh14_w42_8 :  std_logic;
signal bh14_w43_6 :  std_logic;
signal bh14_w44_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid254_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid254_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid254_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid254_Out0_copy255 :  std_logic_vector(2 downto 0);
signal bh14_w44_8 :  std_logic;
signal bh14_w45_6 :  std_logic;
signal bh14_w46_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid256_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid256_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid256_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid256_Out0_copy257 :  std_logic_vector(2 downto 0);
signal bh14_w46_8 :  std_logic;
signal bh14_w47_6 :  std_logic;
signal bh14_w48_8 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid258_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid258_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid258_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid258_Out0_copy259 :  std_logic_vector(2 downto 0);
signal bh14_w48_9 :  std_logic;
signal bh14_w49_7 :  std_logic;
signal bh14_w50_8 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid260_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid260_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid260_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid260_Out0_copy261 :  std_logic_vector(2 downto 0);
signal bh14_w50_9 :  std_logic;
signal bh14_w51_9 :  std_logic;
signal bh14_w52_8 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid262_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid262_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid262_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid262_Out0_copy263 :  std_logic_vector(2 downto 0);
signal bh14_w51_10 :  std_logic;
signal bh14_w52_9 :  std_logic;
signal bh14_w53_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid264_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid264_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid264_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid264_Out0_copy265 :  std_logic_vector(2 downto 0);
signal bh14_w53_10 :  std_logic;
signal bh14_w54_9 :  std_logic;
signal bh14_w55_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid266_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid266_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid266_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid266_Out0_copy267 :  std_logic_vector(2 downto 0);
signal bh14_w55_10 :  std_logic;
signal bh14_w56_9 :  std_logic;
signal bh14_w57_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid268_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid268_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid268_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid268_Out0_copy269 :  std_logic_vector(2 downto 0);
signal bh14_w57_10 :  std_logic;
signal bh14_w58_9 :  std_logic;
signal bh14_w59_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid270_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid270_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid270_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid270_Out0_copy271 :  std_logic_vector(2 downto 0);
signal bh14_w59_10 :  std_logic;
signal bh14_w60_9 :  std_logic;
signal bh14_w61_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid272_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid272_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid272_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid272_Out0_copy273 :  std_logic_vector(2 downto 0);
signal bh14_w61_10 :  std_logic;
signal bh14_w62_9 :  std_logic;
signal bh14_w63_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid274_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid274_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid274_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid274_Out0_copy275 :  std_logic_vector(2 downto 0);
signal bh14_w63_10 :  std_logic;
signal bh14_w64_9 :  std_logic;
signal bh14_w65_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid276_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid276_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid276_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid276_Out0_copy277 :  std_logic_vector(2 downto 0);
signal bh14_w65_10 :  std_logic;
signal bh14_w66_9 :  std_logic;
signal bh14_w67_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid278_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid278_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid278_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid278_Out0_copy279 :  std_logic_vector(2 downto 0);
signal bh14_w67_10 :  std_logic;
signal bh14_w68_9 :  std_logic;
signal bh14_w69_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid280_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid280_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid280_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid280_Out0_copy281 :  std_logic_vector(2 downto 0);
signal bh14_w69_10 :  std_logic;
signal bh14_w70_9 :  std_logic;
signal bh14_w71_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid282_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid282_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid282_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid282_Out0_copy283 :  std_logic_vector(2 downto 0);
signal bh14_w71_10 :  std_logic;
signal bh14_w72_9 :  std_logic;
signal bh14_w73_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid284_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid284_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid284_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid284_Out0_copy285 :  std_logic_vector(2 downto 0);
signal bh14_w73_10 :  std_logic;
signal bh14_w74_9 :  std_logic;
signal bh14_w75_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid286_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid286_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid286_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid286_Out0_copy287 :  std_logic_vector(2 downto 0);
signal bh14_w75_10 :  std_logic;
signal bh14_w76_9 :  std_logic;
signal bh14_w77_10 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid288_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid288_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid288_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid288_Out0_copy289 :  std_logic_vector(2 downto 0);
signal bh14_w77_11 :  std_logic;
signal bh14_w78_9 :  std_logic;
signal bh14_w79_9 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid290_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid290_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid290_Out0_copy291 :  std_logic_vector(1 downto 0);
signal bh14_w78_10 :  std_logic;
signal bh14_w79_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid292_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid292_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid292_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid292_Out0_copy293 :  std_logic_vector(2 downto 0);
signal bh14_w79_11 :  std_logic;
signal bh14_w80_9 :  std_logic;
signal bh14_w81_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid294_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid294_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid294_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid294_Out0_copy295 :  std_logic_vector(2 downto 0);
signal bh14_w81_10 :  std_logic;
signal bh14_w82_9 :  std_logic;
signal bh14_w83_9 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid296_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid296_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid296_Out0_copy297 :  std_logic_vector(1 downto 0);
signal bh14_w83_10 :  std_logic;
signal bh14_w84_8 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid298_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid298_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid298_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid298_Out0_copy299 :  std_logic_vector(2 downto 0);
signal bh14_w84_9 :  std_logic;
signal bh14_w85_8 :  std_logic;
signal bh14_w86_8 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid300_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid300_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid300_Out0_copy301 :  std_logic_vector(1 downto 0);
signal bh14_w85_9 :  std_logic;
signal bh14_w86_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid302_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid302_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid302_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid302_Out0_copy303 :  std_logic_vector(2 downto 0);
signal bh14_w86_10 :  std_logic;
signal bh14_w87_8 :  std_logic;
signal bh14_w88_8 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid304_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid304_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid304_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid304_Out0_copy305 :  std_logic_vector(2 downto 0);
signal bh14_w88_9 :  std_logic;
signal bh14_w89_8 :  std_logic;
signal bh14_w90_8 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid306_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid306_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid306_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid306_Out0_copy307 :  std_logic_vector(2 downto 0);
signal bh14_w90_9 :  std_logic;
signal bh14_w91_8 :  std_logic;
signal bh14_w92_8 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid308_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid308_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid308_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid308_Out0_copy309 :  std_logic_vector(2 downto 0);
signal bh14_w92_9 :  std_logic;
signal bh14_w93_8 :  std_logic;
signal bh14_w94_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid310_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid310_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid310_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid310_Out0_copy311 :  std_logic_vector(2 downto 0);
signal bh14_w94_8 :  std_logic;
signal bh14_w95_7 :  std_logic;
signal bh14_w96_6 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid312_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid312_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid312_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid312_Out0_copy313 :  std_logic_vector(2 downto 0);
signal bh14_w95_8 :  std_logic;
signal bh14_w96_7 :  std_logic;
signal bh14_w97_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid314_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid314_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid314_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid314_Out0_copy315 :  std_logic_vector(2 downto 0);
signal bh14_w97_8 :  std_logic;
signal bh14_w98_6 :  std_logic;
signal bh14_w99_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid316_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid316_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid316_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid316_Out0_copy317 :  std_logic_vector(2 downto 0);
signal bh14_w99_8 :  std_logic;
signal bh14_w100_6 :  std_logic;
signal bh14_w101_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid318_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid318_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid318_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid318_Out0_copy319 :  std_logic_vector(2 downto 0);
signal bh14_w101_8 :  std_logic;
signal bh14_w102_6 :  std_logic;
signal bh14_w103_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid320_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid320_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid320_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid320_Out0_copy321 :  std_logic_vector(2 downto 0);
signal bh14_w103_8 :  std_logic;
signal bh14_w104_6 :  std_logic;
signal bh14_w105_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid322_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid322_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid322_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid322_Out0_copy323 :  std_logic_vector(2 downto 0);
signal bh14_w105_8 :  std_logic;
signal bh14_w106_6 :  std_logic;
signal bh14_w107_7 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid324_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid324_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid324_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid324_Out0_copy325 :  std_logic_vector(2 downto 0);
signal bh14_w107_8 :  std_logic;
signal bh14_w108_5 :  std_logic;
signal bh14_w109_6 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid326_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid326_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid326_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid326_Out0_copy327 :  std_logic_vector(2 downto 0);
signal bh14_w109_7 :  std_logic;
signal bh14_w110_4 :  std_logic;
signal bh14_w111_4 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid328_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid328_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid328_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid328_Out0_copy329 :  std_logic_vector(2 downto 0);
signal bh14_w111_5 :  std_logic;
signal bh14_w112_3 :  std_logic;
signal bh14_w113_4 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid330_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid330_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid330_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid330_Out0_copy331 :  std_logic_vector(2 downto 0);
signal bh14_w113_5 :  std_logic;
signal bh14_w114_3 :  std_logic;
signal bh14_w115_4 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid332_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid332_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid332_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid332_Out0_copy333 :  std_logic_vector(2 downto 0);
signal bh14_w115_5 :  std_logic;
signal bh14_w116_3 :  std_logic;
signal bh14_w117_4 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid334_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid334_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid334_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid334_Out0_copy335 :  std_logic_vector(2 downto 0);
signal bh14_w117_5 :  std_logic;
signal bh14_w118_3 :  std_logic;
signal bh14_w119_4 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid336_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid336_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid336_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid336_Out0_copy337 :  std_logic_vector(2 downto 0);
signal bh14_w119_5 :  std_logic;
signal bh14_w120_3 :  std_logic;
signal bh14_w121_2 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid338_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid338_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid338_Out0_copy339 :  std_logic_vector(1 downto 0);
signal bh14_w121_3 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid340_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid340_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid340_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid340_Out0_copy341 :  std_logic_vector(2 downto 0);
signal bh14_w21_6 :  std_logic;
signal bh14_w22_4 :  std_logic;
signal bh14_w23_6 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid342_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid342_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid342_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid342_Out0_copy343 :  std_logic_vector(2 downto 0);
signal bh14_w23_7 :  std_logic;
signal bh14_w24_6 :  std_logic;
signal bh14_w25_6 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid344_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid344_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid344_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid344_Out0_copy345 :  std_logic_vector(2 downto 0);
signal bh14_w25_7 :  std_logic;
signal bh14_w26_6 :  std_logic;
signal bh14_w27_6 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid346_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid346_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid346_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid346_Out0_copy347 :  std_logic_vector(2 downto 0);
signal bh14_w27_7 :  std_logic;
signal bh14_w28_6 :  std_logic;
signal bh14_w29_6 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid348_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid348_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid348_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid348_Out0_copy349 :  std_logic_vector(2 downto 0);
signal bh14_w29_7 :  std_logic;
signal bh14_w30_6 :  std_logic;
signal bh14_w31_6 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid350_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid350_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid350_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid350_Out0_copy351 :  std_logic_vector(2 downto 0);
signal bh14_w31_7 :  std_logic;
signal bh14_w32_6 :  std_logic;
signal bh14_w33_6 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid352_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid352_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid352_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid352_Out0_copy353 :  std_logic_vector(2 downto 0);
signal bh14_w33_7 :  std_logic;
signal bh14_w34_7 :  std_logic;
signal bh14_w35_8 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid354_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid354_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid354_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid354_Out0_copy355 :  std_logic_vector(2 downto 0);
signal bh14_w35_9 :  std_logic;
signal bh14_w36_9 :  std_logic;
signal bh14_w37_7 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid356_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid356_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid356_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid356_Out0_copy357 :  std_logic_vector(2 downto 0);
signal bh14_w38_9 :  std_logic;
signal bh14_w39_7 :  std_logic;
signal bh14_w40_9 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid358_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid358_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid358_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid358_Out0_copy359 :  std_logic_vector(2 downto 0);
signal bh14_w40_10 :  std_logic;
signal bh14_w41_7 :  std_logic;
signal bh14_w42_9 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid360_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid360_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid360_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid360_Out0_copy361 :  std_logic_vector(2 downto 0);
signal bh14_w42_10 :  std_logic;
signal bh14_w43_7 :  std_logic;
signal bh14_w44_9 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid362_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid362_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid362_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid362_Out0_copy363 :  std_logic_vector(2 downto 0);
signal bh14_w44_10 :  std_logic;
signal bh14_w45_7 :  std_logic;
signal bh14_w46_9 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid364_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid364_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid364_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid364_Out0_copy365 :  std_logic_vector(2 downto 0);
signal bh14_w46_10 :  std_logic;
signal bh14_w47_7 :  std_logic;
signal bh14_w48_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid366_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid366_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid366_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid366_Out0_copy367 :  std_logic_vector(2 downto 0);
signal bh14_w48_11 :  std_logic;
signal bh14_w49_8 :  std_logic;
signal bh14_w50_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid368_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid368_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid368_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid368_Out0_copy369 :  std_logic_vector(2 downto 0);
signal bh14_w50_11 :  std_logic;
signal bh14_w51_11 :  std_logic;
signal bh14_w52_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid370_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid370_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid370_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid370_Out0_copy371 :  std_logic_vector(2 downto 0);
signal bh14_w52_11 :  std_logic;
signal bh14_w53_11 :  std_logic;
signal bh14_w54_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid372_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid372_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid372_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid372_Out0_copy373 :  std_logic_vector(2 downto 0);
signal bh14_w54_11 :  std_logic;
signal bh14_w55_11 :  std_logic;
signal bh14_w56_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid374_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid374_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid374_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid374_Out0_copy375 :  std_logic_vector(2 downto 0);
signal bh14_w56_11 :  std_logic;
signal bh14_w57_11 :  std_logic;
signal bh14_w58_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid376_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid376_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid376_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid376_Out0_copy377 :  std_logic_vector(2 downto 0);
signal bh14_w58_11 :  std_logic;
signal bh14_w59_11 :  std_logic;
signal bh14_w60_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid378_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid378_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid378_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid378_Out0_copy379 :  std_logic_vector(2 downto 0);
signal bh14_w60_11 :  std_logic;
signal bh14_w61_11 :  std_logic;
signal bh14_w62_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid380_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid380_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid380_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid380_Out0_copy381 :  std_logic_vector(2 downto 0);
signal bh14_w62_11 :  std_logic;
signal bh14_w63_11 :  std_logic;
signal bh14_w64_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid382_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid382_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid382_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid382_Out0_copy383 :  std_logic_vector(2 downto 0);
signal bh14_w64_11 :  std_logic;
signal bh14_w65_11 :  std_logic;
signal bh14_w66_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid384_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid384_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid384_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid384_Out0_copy385 :  std_logic_vector(2 downto 0);
signal bh14_w66_11 :  std_logic;
signal bh14_w67_11 :  std_logic;
signal bh14_w68_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid386_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid386_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid386_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid386_Out0_copy387 :  std_logic_vector(2 downto 0);
signal bh14_w68_11 :  std_logic;
signal bh14_w69_11 :  std_logic;
signal bh14_w70_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid388_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid388_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid388_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid388_Out0_copy389 :  std_logic_vector(2 downto 0);
signal bh14_w70_11 :  std_logic;
signal bh14_w71_11 :  std_logic;
signal bh14_w72_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid390_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid390_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid390_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid390_Out0_copy391 :  std_logic_vector(2 downto 0);
signal bh14_w72_11 :  std_logic;
signal bh14_w73_11 :  std_logic;
signal bh14_w74_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid392_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid392_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid392_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid392_Out0_copy393 :  std_logic_vector(2 downto 0);
signal bh14_w74_11 :  std_logic;
signal bh14_w75_11 :  std_logic;
signal bh14_w76_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid394_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid394_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid394_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid394_Out0_copy395 :  std_logic_vector(2 downto 0);
signal bh14_w76_11 :  std_logic;
signal bh14_w77_12 :  std_logic;
signal bh14_w78_11 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid396_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid396_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid396_Out0_copy397 :  std_logic_vector(1 downto 0);
signal bh14_w78_12 :  std_logic;
signal bh14_w79_12 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid398_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid398_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid398_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid398_Out0_copy399 :  std_logic_vector(2 downto 0);
signal bh14_w79_13 :  std_logic;
signal bh14_w80_10 :  std_logic;
signal bh14_w81_11 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid400_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid400_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid400_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid400_Out0_copy401 :  std_logic_vector(2 downto 0);
signal bh14_w81_12 :  std_logic;
signal bh14_w82_10 :  std_logic;
signal bh14_w83_11 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid402_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid402_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid402_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid402_Out0_copy403 :  std_logic_vector(2 downto 0);
signal bh14_w83_12 :  std_logic;
signal bh14_w84_10 :  std_logic;
signal bh14_w85_10 :  std_logic;
signal Compressor_3_2_F50_uid49_bh14_uid404_In0 :  std_logic_vector(2 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid404_Out0 :  std_logic_vector(1 downto 0);
signal Compressor_3_2_F50_uid49_bh14_uid404_Out0_copy405 :  std_logic_vector(1 downto 0);
signal bh14_w85_11 :  std_logic;
signal bh14_w86_11 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid406_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid406_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid406_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid406_Out0_copy407 :  std_logic_vector(2 downto 0);
signal bh14_w86_12 :  std_logic;
signal bh14_w87_9 :  std_logic;
signal bh14_w88_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid408_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid408_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid408_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid408_Out0_copy409 :  std_logic_vector(2 downto 0);
signal bh14_w88_11 :  std_logic;
signal bh14_w89_9 :  std_logic;
signal bh14_w90_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid410_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid410_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid410_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid410_Out0_copy411 :  std_logic_vector(2 downto 0);
signal bh14_w90_11 :  std_logic;
signal bh14_w91_9 :  std_logic;
signal bh14_w92_10 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid412_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid412_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid412_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid412_Out0_copy413 :  std_logic_vector(2 downto 0);
signal bh14_w92_11 :  std_logic;
signal bh14_w93_9 :  std_logic;
signal bh14_w94_9 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid414_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid414_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid414_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid414_Out0_copy415 :  std_logic_vector(2 downto 0);
signal bh14_w94_10 :  std_logic;
signal bh14_w95_9 :  std_logic;
signal bh14_w96_8 :  std_logic;
signal Compressor_23_3_F50_uid41_bh14_uid416_In0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid416_In1 :  std_logic_vector(1 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid416_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_23_3_F50_uid41_bh14_uid416_Out0_copy417 :  std_logic_vector(2 downto 0);
signal bh14_w96_9 :  std_logic;
signal bh14_w97_9 :  std_logic;
signal bh14_w98_7 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid418_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid418_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid418_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid418_Out0_copy419 :  std_logic_vector(2 downto 0);
signal bh14_w99_9 :  std_logic;
signal bh14_w100_7 :  std_logic;
signal bh14_w101_9 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid420_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid420_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid420_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid420_Out0_copy421 :  std_logic_vector(2 downto 0);
signal bh14_w101_10 :  std_logic;
signal bh14_w102_7 :  std_logic;
signal bh14_w103_9 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid422_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid422_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid422_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid422_Out0_copy423 :  std_logic_vector(2 downto 0);
signal bh14_w103_10 :  std_logic;
signal bh14_w104_7 :  std_logic;
signal bh14_w105_9 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid424_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid424_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid424_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid424_Out0_copy425 :  std_logic_vector(2 downto 0);
signal bh14_w105_10 :  std_logic;
signal bh14_w106_7 :  std_logic;
signal bh14_w107_9 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid426_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid426_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid426_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid426_Out0_copy427 :  std_logic_vector(2 downto 0);
signal bh14_w107_10 :  std_logic;
signal bh14_w108_6 :  std_logic;
signal bh14_w109_8 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid428_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid428_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid428_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid428_Out0_copy429 :  std_logic_vector(2 downto 0);
signal bh14_w109_9 :  std_logic;
signal bh14_w110_5 :  std_logic;
signal bh14_w111_6 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid430_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid430_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid430_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid430_Out0_copy431 :  std_logic_vector(2 downto 0);
signal bh14_w111_7 :  std_logic;
signal bh14_w112_4 :  std_logic;
signal bh14_w113_6 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid432_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid432_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid432_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid432_Out0_copy433 :  std_logic_vector(2 downto 0);
signal bh14_w113_7 :  std_logic;
signal bh14_w114_4 :  std_logic;
signal bh14_w115_6 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid434_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid434_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid434_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid434_Out0_copy435 :  std_logic_vector(2 downto 0);
signal bh14_w115_7 :  std_logic;
signal bh14_w116_4 :  std_logic;
signal bh14_w117_6 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid436_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid436_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid436_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid436_Out0_copy437 :  std_logic_vector(2 downto 0);
signal bh14_w117_7 :  std_logic;
signal bh14_w118_4 :  std_logic;
signal bh14_w119_6 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid438_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid438_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid438_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid438_Out0_copy439 :  std_logic_vector(2 downto 0);
signal bh14_w119_7 :  std_logic;
signal bh14_w120_4 :  std_logic;
signal bh14_w121_4 :  std_logic;
signal Compressor_14_3_F50_uid63_bh14_uid440_In0 :  std_logic_vector(3 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid440_In1 :  std_logic_vector(0 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid440_Out0 :  std_logic_vector(2 downto 0);
signal Compressor_14_3_F50_uid63_bh14_uid440_Out0_copy441 :  std_logic_vector(2 downto 0);
signal bh14_w121_5 :  std_logic;
signal tmp_bitheapResult_bh14_22 :  std_logic_vector(22 downto 0);
signal bitheapFinalAdd_bh14_In0 :  std_logic_vector(99 downto 0);
signal bitheapFinalAdd_bh14_In1 :  std_logic_vector(99 downto 0);
signal bitheapFinalAdd_bh14_Cin :  std_logic;
signal bitheapFinalAdd_bh14_Out :  std_logic_vector(99 downto 0);
signal bitheapResult_bh14 :  std_logic_vector(121 downto 0);
begin
   XX_m13 <= X ;
   YY_m13 <= Y ;
   tile_0_X <= X(16 downto 0);
   tile_0_Y <= Y(23 downto 0);
   tile_0_mult: DSPBlock_17x24_F50_uid16
      port map ( clk  => clk,
                 X => tile_0_X,
                 Y => tile_0_Y,
                 R => tile_0_output);

   tile_0_filtered_output <= unsigned(tile_0_output(40 downto 0));
   bh14_w0_0 <= tile_0_filtered_output(0);
   bh14_w1_0 <= tile_0_filtered_output(1);
   bh14_w2_0 <= tile_0_filtered_output(2);
   bh14_w3_0 <= tile_0_filtered_output(3);
   bh14_w4_0 <= tile_0_filtered_output(4);
   bh14_w5_0 <= tile_0_filtered_output(5);
   bh14_w6_0 <= tile_0_filtered_output(6);
   bh14_w7_0 <= tile_0_filtered_output(7);
   bh14_w8_0 <= tile_0_filtered_output(8);
   bh14_w9_0 <= tile_0_filtered_output(9);
   bh14_w10_0 <= tile_0_filtered_output(10);
   bh14_w11_0 <= tile_0_filtered_output(11);
   bh14_w12_0 <= tile_0_filtered_output(12);
   bh14_w13_0 <= tile_0_filtered_output(13);
   bh14_w14_0 <= tile_0_filtered_output(14);
   bh14_w15_0 <= tile_0_filtered_output(15);
   bh14_w16_0 <= tile_0_filtered_output(16);
   bh14_w17_0 <= tile_0_filtered_output(17);
   bh14_w18_0 <= tile_0_filtered_output(18);
   bh14_w19_0 <= tile_0_filtered_output(19);
   bh14_w20_0 <= tile_0_filtered_output(20);
   bh14_w21_0 <= tile_0_filtered_output(21);
   bh14_w22_0 <= tile_0_filtered_output(22);
   bh14_w23_0 <= tile_0_filtered_output(23);
   bh14_w24_0 <= tile_0_filtered_output(24);
   bh14_w25_0 <= tile_0_filtered_output(25);
   bh14_w26_0 <= tile_0_filtered_output(26);
   bh14_w27_0 <= tile_0_filtered_output(27);
   bh14_w28_0 <= tile_0_filtered_output(28);
   bh14_w29_0 <= tile_0_filtered_output(29);
   bh14_w30_0 <= tile_0_filtered_output(30);
   bh14_w31_0 <= tile_0_filtered_output(31);
   bh14_w32_0 <= tile_0_filtered_output(32);
   bh14_w33_0 <= tile_0_filtered_output(33);
   bh14_w34_0 <= tile_0_filtered_output(34);
   bh14_w35_0 <= tile_0_filtered_output(35);
   bh14_w36_0 <= tile_0_filtered_output(36);
   bh14_w37_0 <= tile_0_filtered_output(37);
   bh14_w38_0 <= tile_0_filtered_output(38);
   bh14_w39_0 <= tile_0_filtered_output(39);
   bh14_w40_0 <= tile_0_filtered_output(40);
   tile_1_X <= X(33 downto 17);
   tile_1_Y <= Y(23 downto 0);
   tile_1_mult: DSPBlock_17x24_F50_uid18
      port map ( clk  => clk,
                 X => tile_1_X,
                 Y => tile_1_Y,
                 R => tile_1_output);

   tile_1_filtered_output <= unsigned(tile_1_output(40 downto 0));
   bh14_w17_1 <= tile_1_filtered_output(0);
   bh14_w18_1 <= tile_1_filtered_output(1);
   bh14_w19_1 <= tile_1_filtered_output(2);
   bh14_w20_1 <= tile_1_filtered_output(3);
   bh14_w21_1 <= tile_1_filtered_output(4);
   bh14_w22_1 <= tile_1_filtered_output(5);
   bh14_w23_1 <= tile_1_filtered_output(6);
   bh14_w24_1 <= tile_1_filtered_output(7);
   bh14_w25_1 <= tile_1_filtered_output(8);
   bh14_w26_1 <= tile_1_filtered_output(9);
   bh14_w27_1 <= tile_1_filtered_output(10);
   bh14_w28_1 <= tile_1_filtered_output(11);
   bh14_w29_1 <= tile_1_filtered_output(12);
   bh14_w30_1 <= tile_1_filtered_output(13);
   bh14_w31_1 <= tile_1_filtered_output(14);
   bh14_w32_1 <= tile_1_filtered_output(15);
   bh14_w33_1 <= tile_1_filtered_output(16);
   bh14_w34_1 <= tile_1_filtered_output(17);
   bh14_w35_1 <= tile_1_filtered_output(18);
   bh14_w36_1 <= tile_1_filtered_output(19);
   bh14_w37_1 <= tile_1_filtered_output(20);
   bh14_w38_1 <= tile_1_filtered_output(21);
   bh14_w39_1 <= tile_1_filtered_output(22);
   bh14_w40_1 <= tile_1_filtered_output(23);
   bh14_w41_0 <= tile_1_filtered_output(24);
   bh14_w42_0 <= tile_1_filtered_output(25);
   bh14_w43_0 <= tile_1_filtered_output(26);
   bh14_w44_0 <= tile_1_filtered_output(27);
   bh14_w45_0 <= tile_1_filtered_output(28);
   bh14_w46_0 <= tile_1_filtered_output(29);
   bh14_w47_0 <= tile_1_filtered_output(30);
   bh14_w48_0 <= tile_1_filtered_output(31);
   bh14_w49_0 <= tile_1_filtered_output(32);
   bh14_w50_0 <= tile_1_filtered_output(33);
   bh14_w51_0 <= tile_1_filtered_output(34);
   bh14_w52_0 <= tile_1_filtered_output(35);
   bh14_w53_0 <= tile_1_filtered_output(36);
   bh14_w54_0 <= tile_1_filtered_output(37);
   bh14_w55_0 <= tile_1_filtered_output(38);
   bh14_w56_0 <= tile_1_filtered_output(39);
   bh14_w57_0 <= tile_1_filtered_output(40);
   tile_2_X <= X(50 downto 34);
   tile_2_Y <= Y(23 downto 0);
   tile_2_mult: DSPBlock_17x24_F50_uid20
      port map ( clk  => clk,
                 X => tile_2_X,
                 Y => tile_2_Y,
                 R => tile_2_output);

   tile_2_filtered_output <= unsigned(tile_2_output(40 downto 0));
   bh14_w34_2 <= tile_2_filtered_output(0);
   bh14_w35_2 <= tile_2_filtered_output(1);
   bh14_w36_2 <= tile_2_filtered_output(2);
   bh14_w37_2 <= tile_2_filtered_output(3);
   bh14_w38_2 <= tile_2_filtered_output(4);
   bh14_w39_2 <= tile_2_filtered_output(5);
   bh14_w40_2 <= tile_2_filtered_output(6);
   bh14_w41_1 <= tile_2_filtered_output(7);
   bh14_w42_1 <= tile_2_filtered_output(8);
   bh14_w43_1 <= tile_2_filtered_output(9);
   bh14_w44_1 <= tile_2_filtered_output(10);
   bh14_w45_1 <= tile_2_filtered_output(11);
   bh14_w46_1 <= tile_2_filtered_output(12);
   bh14_w47_1 <= tile_2_filtered_output(13);
   bh14_w48_1 <= tile_2_filtered_output(14);
   bh14_w49_1 <= tile_2_filtered_output(15);
   bh14_w50_1 <= tile_2_filtered_output(16);
   bh14_w51_1 <= tile_2_filtered_output(17);
   bh14_w52_1 <= tile_2_filtered_output(18);
   bh14_w53_1 <= tile_2_filtered_output(19);
   bh14_w54_1 <= tile_2_filtered_output(20);
   bh14_w55_1 <= tile_2_filtered_output(21);
   bh14_w56_1 <= tile_2_filtered_output(22);
   bh14_w57_1 <= tile_2_filtered_output(23);
   bh14_w58_0 <= tile_2_filtered_output(24);
   bh14_w59_0 <= tile_2_filtered_output(25);
   bh14_w60_0 <= tile_2_filtered_output(26);
   bh14_w61_0 <= tile_2_filtered_output(27);
   bh14_w62_0 <= tile_2_filtered_output(28);
   bh14_w63_0 <= tile_2_filtered_output(29);
   bh14_w64_0 <= tile_2_filtered_output(30);
   bh14_w65_0 <= tile_2_filtered_output(31);
   bh14_w66_0 <= tile_2_filtered_output(32);
   bh14_w67_0 <= tile_2_filtered_output(33);
   bh14_w68_0 <= tile_2_filtered_output(34);
   bh14_w69_0 <= tile_2_filtered_output(35);
   bh14_w70_0 <= tile_2_filtered_output(36);
   bh14_w71_0 <= tile_2_filtered_output(37);
   bh14_w72_0 <= tile_2_filtered_output(38);
   bh14_w73_0 <= tile_2_filtered_output(39);
   bh14_w74_0 <= tile_2_filtered_output(40);
   tile_3_X <= X(60 downto 51);
   tile_3_Y <= Y(23 downto 0);
   tile_3_mult: DSPBlock_10x24_F50_uid22
      port map ( clk  => clk,
                 X => tile_3_X,
                 Y => tile_3_Y,
                 R => tile_3_output);

   tile_3_filtered_output <= signed(tile_3_output(33 downto 0));
   bh14_w51_2 <= tile_3_filtered_output(0);
   bh14_w52_2 <= tile_3_filtered_output(1);
   bh14_w53_2 <= tile_3_filtered_output(2);
   bh14_w54_2 <= tile_3_filtered_output(3);
   bh14_w55_2 <= tile_3_filtered_output(4);
   bh14_w56_2 <= tile_3_filtered_output(5);
   bh14_w57_2 <= tile_3_filtered_output(6);
   bh14_w58_1 <= tile_3_filtered_output(7);
   bh14_w59_1 <= tile_3_filtered_output(8);
   bh14_w60_1 <= tile_3_filtered_output(9);
   bh14_w61_1 <= tile_3_filtered_output(10);
   bh14_w62_1 <= tile_3_filtered_output(11);
   bh14_w63_1 <= tile_3_filtered_output(12);
   bh14_w64_1 <= tile_3_filtered_output(13);
   bh14_w65_1 <= tile_3_filtered_output(14);
   bh14_w66_1 <= tile_3_filtered_output(15);
   bh14_w67_1 <= tile_3_filtered_output(16);
   bh14_w68_1 <= tile_3_filtered_output(17);
   bh14_w69_1 <= tile_3_filtered_output(18);
   bh14_w70_1 <= tile_3_filtered_output(19);
   bh14_w71_1 <= tile_3_filtered_output(20);
   bh14_w72_1 <= tile_3_filtered_output(21);
   bh14_w73_1 <= tile_3_filtered_output(22);
   bh14_w74_1 <= tile_3_filtered_output(23);
   bh14_w75_0 <= tile_3_filtered_output(24);
   bh14_w76_0 <= tile_3_filtered_output(25);
   bh14_w77_0 <= tile_3_filtered_output(26);
   bh14_w78_0 <= tile_3_filtered_output(27);
   bh14_w79_0 <= tile_3_filtered_output(28);
   bh14_w80_0 <= tile_3_filtered_output(29);
   bh14_w81_0 <= tile_3_filtered_output(30);
   bh14_w82_0 <= tile_3_filtered_output(31);
   bh14_w83_0 <= tile_3_filtered_output(32);
   bh14_w84_0 <= not tile_3_filtered_output(33);
   tile_4_X <= X(16 downto 0);
   tile_4_Y <= Y(47 downto 24);
   tile_4_mult: DSPBlock_17x24_F50_uid24
      port map ( clk  => clk,
                 X => tile_4_X,
                 Y => tile_4_Y,
                 R => tile_4_output);

   tile_4_filtered_output <= unsigned(tile_4_output(40 downto 0));
   bh14_w24_2 <= tile_4_filtered_output(0);
   bh14_w25_2 <= tile_4_filtered_output(1);
   bh14_w26_2 <= tile_4_filtered_output(2);
   bh14_w27_2 <= tile_4_filtered_output(3);
   bh14_w28_2 <= tile_4_filtered_output(4);
   bh14_w29_2 <= tile_4_filtered_output(5);
   bh14_w30_2 <= tile_4_filtered_output(6);
   bh14_w31_2 <= tile_4_filtered_output(7);
   bh14_w32_2 <= tile_4_filtered_output(8);
   bh14_w33_2 <= tile_4_filtered_output(9);
   bh14_w34_3 <= tile_4_filtered_output(10);
   bh14_w35_3 <= tile_4_filtered_output(11);
   bh14_w36_3 <= tile_4_filtered_output(12);
   bh14_w37_3 <= tile_4_filtered_output(13);
   bh14_w38_3 <= tile_4_filtered_output(14);
   bh14_w39_3 <= tile_4_filtered_output(15);
   bh14_w40_3 <= tile_4_filtered_output(16);
   bh14_w41_2 <= tile_4_filtered_output(17);
   bh14_w42_2 <= tile_4_filtered_output(18);
   bh14_w43_2 <= tile_4_filtered_output(19);
   bh14_w44_2 <= tile_4_filtered_output(20);
   bh14_w45_2 <= tile_4_filtered_output(21);
   bh14_w46_2 <= tile_4_filtered_output(22);
   bh14_w47_2 <= tile_4_filtered_output(23);
   bh14_w48_2 <= tile_4_filtered_output(24);
   bh14_w49_2 <= tile_4_filtered_output(25);
   bh14_w50_2 <= tile_4_filtered_output(26);
   bh14_w51_3 <= tile_4_filtered_output(27);
   bh14_w52_3 <= tile_4_filtered_output(28);
   bh14_w53_3 <= tile_4_filtered_output(29);
   bh14_w54_3 <= tile_4_filtered_output(30);
   bh14_w55_3 <= tile_4_filtered_output(31);
   bh14_w56_3 <= tile_4_filtered_output(32);
   bh14_w57_3 <= tile_4_filtered_output(33);
   bh14_w58_2 <= tile_4_filtered_output(34);
   bh14_w59_2 <= tile_4_filtered_output(35);
   bh14_w60_2 <= tile_4_filtered_output(36);
   bh14_w61_2 <= tile_4_filtered_output(37);
   bh14_w62_2 <= tile_4_filtered_output(38);
   bh14_w63_2 <= tile_4_filtered_output(39);
   bh14_w64_2 <= tile_4_filtered_output(40);
   tile_5_X <= X(33 downto 17);
   tile_5_Y <= Y(47 downto 24);
   tile_5_mult: DSPBlock_17x24_F50_uid26
      port map ( clk  => clk,
                 X => tile_5_X,
                 Y => tile_5_Y,
                 R => tile_5_output);

   tile_5_filtered_output <= unsigned(tile_5_output(40 downto 0));
   bh14_w41_3 <= tile_5_filtered_output(0);
   bh14_w42_3 <= tile_5_filtered_output(1);
   bh14_w43_3 <= tile_5_filtered_output(2);
   bh14_w44_3 <= tile_5_filtered_output(3);
   bh14_w45_3 <= tile_5_filtered_output(4);
   bh14_w46_3 <= tile_5_filtered_output(5);
   bh14_w47_3 <= tile_5_filtered_output(6);
   bh14_w48_3 <= tile_5_filtered_output(7);
   bh14_w49_3 <= tile_5_filtered_output(8);
   bh14_w50_3 <= tile_5_filtered_output(9);
   bh14_w51_4 <= tile_5_filtered_output(10);
   bh14_w52_4 <= tile_5_filtered_output(11);
   bh14_w53_4 <= tile_5_filtered_output(12);
   bh14_w54_4 <= tile_5_filtered_output(13);
   bh14_w55_4 <= tile_5_filtered_output(14);
   bh14_w56_4 <= tile_5_filtered_output(15);
   bh14_w57_4 <= tile_5_filtered_output(16);
   bh14_w58_3 <= tile_5_filtered_output(17);
   bh14_w59_3 <= tile_5_filtered_output(18);
   bh14_w60_3 <= tile_5_filtered_output(19);
   bh14_w61_3 <= tile_5_filtered_output(20);
   bh14_w62_3 <= tile_5_filtered_output(21);
   bh14_w63_3 <= tile_5_filtered_output(22);
   bh14_w64_3 <= tile_5_filtered_output(23);
   bh14_w65_2 <= tile_5_filtered_output(24);
   bh14_w66_2 <= tile_5_filtered_output(25);
   bh14_w67_2 <= tile_5_filtered_output(26);
   bh14_w68_2 <= tile_5_filtered_output(27);
   bh14_w69_2 <= tile_5_filtered_output(28);
   bh14_w70_2 <= tile_5_filtered_output(29);
   bh14_w71_2 <= tile_5_filtered_output(30);
   bh14_w72_2 <= tile_5_filtered_output(31);
   bh14_w73_2 <= tile_5_filtered_output(32);
   bh14_w74_2 <= tile_5_filtered_output(33);
   bh14_w75_1 <= tile_5_filtered_output(34);
   bh14_w76_1 <= tile_5_filtered_output(35);
   bh14_w77_1 <= tile_5_filtered_output(36);
   bh14_w78_1 <= tile_5_filtered_output(37);
   bh14_w79_1 <= tile_5_filtered_output(38);
   bh14_w80_1 <= tile_5_filtered_output(39);
   bh14_w81_1 <= tile_5_filtered_output(40);
   tile_6_X <= X(50 downto 34);
   tile_6_Y <= Y(47 downto 24);
   tile_6_mult: DSPBlock_17x24_F50_uid28
      port map ( clk  => clk,
                 X => tile_6_X,
                 Y => tile_6_Y,
                 R => tile_6_output);

   tile_6_filtered_output <= unsigned(tile_6_output(40 downto 0));
   bh14_w58_4 <= tile_6_filtered_output(0);
   bh14_w59_4 <= tile_6_filtered_output(1);
   bh14_w60_4 <= tile_6_filtered_output(2);
   bh14_w61_4 <= tile_6_filtered_output(3);
   bh14_w62_4 <= tile_6_filtered_output(4);
   bh14_w63_4 <= tile_6_filtered_output(5);
   bh14_w64_4 <= tile_6_filtered_output(6);
   bh14_w65_3 <= tile_6_filtered_output(7);
   bh14_w66_3 <= tile_6_filtered_output(8);
   bh14_w67_3 <= tile_6_filtered_output(9);
   bh14_w68_3 <= tile_6_filtered_output(10);
   bh14_w69_3 <= tile_6_filtered_output(11);
   bh14_w70_3 <= tile_6_filtered_output(12);
   bh14_w71_3 <= tile_6_filtered_output(13);
   bh14_w72_3 <= tile_6_filtered_output(14);
   bh14_w73_3 <= tile_6_filtered_output(15);
   bh14_w74_3 <= tile_6_filtered_output(16);
   bh14_w75_2 <= tile_6_filtered_output(17);
   bh14_w76_2 <= tile_6_filtered_output(18);
   bh14_w77_2 <= tile_6_filtered_output(19);
   bh14_w78_2 <= tile_6_filtered_output(20);
   bh14_w79_2 <= tile_6_filtered_output(21);
   bh14_w80_2 <= tile_6_filtered_output(22);
   bh14_w81_2 <= tile_6_filtered_output(23);
   bh14_w82_1 <= tile_6_filtered_output(24);
   bh14_w83_1 <= tile_6_filtered_output(25);
   bh14_w84_1 <= tile_6_filtered_output(26);
   bh14_w85_0 <= tile_6_filtered_output(27);
   bh14_w86_0 <= tile_6_filtered_output(28);
   bh14_w87_0 <= tile_6_filtered_output(29);
   bh14_w88_0 <= tile_6_filtered_output(30);
   bh14_w89_0 <= tile_6_filtered_output(31);
   bh14_w90_0 <= tile_6_filtered_output(32);
   bh14_w91_0 <= tile_6_filtered_output(33);
   bh14_w92_0 <= tile_6_filtered_output(34);
   bh14_w93_0 <= tile_6_filtered_output(35);
   bh14_w94_0 <= tile_6_filtered_output(36);
   bh14_w95_0 <= tile_6_filtered_output(37);
   bh14_w96_0 <= tile_6_filtered_output(38);
   bh14_w97_0 <= tile_6_filtered_output(39);
   bh14_w98_0 <= tile_6_filtered_output(40);
   tile_7_X <= X(60 downto 51);
   tile_7_Y <= Y(47 downto 24);
   tile_7_mult: DSPBlock_10x24_F50_uid30
      port map ( clk  => clk,
                 X => tile_7_X,
                 Y => tile_7_Y,
                 R => tile_7_output);

   tile_7_filtered_output <= signed(tile_7_output(33 downto 0));
   bh14_w75_3 <= tile_7_filtered_output(0);
   bh14_w76_3 <= tile_7_filtered_output(1);
   bh14_w77_3 <= tile_7_filtered_output(2);
   bh14_w78_3 <= tile_7_filtered_output(3);
   bh14_w79_3 <= tile_7_filtered_output(4);
   bh14_w80_3 <= tile_7_filtered_output(5);
   bh14_w81_3 <= tile_7_filtered_output(6);
   bh14_w82_2 <= tile_7_filtered_output(7);
   bh14_w83_2 <= tile_7_filtered_output(8);
   bh14_w84_2 <= tile_7_filtered_output(9);
   bh14_w85_1 <= tile_7_filtered_output(10);
   bh14_w86_1 <= tile_7_filtered_output(11);
   bh14_w87_1 <= tile_7_filtered_output(12);
   bh14_w88_1 <= tile_7_filtered_output(13);
   bh14_w89_1 <= tile_7_filtered_output(14);
   bh14_w90_1 <= tile_7_filtered_output(15);
   bh14_w91_1 <= tile_7_filtered_output(16);
   bh14_w92_1 <= tile_7_filtered_output(17);
   bh14_w93_1 <= tile_7_filtered_output(18);
   bh14_w94_1 <= tile_7_filtered_output(19);
   bh14_w95_1 <= tile_7_filtered_output(20);
   bh14_w96_1 <= tile_7_filtered_output(21);
   bh14_w97_1 <= tile_7_filtered_output(22);
   bh14_w98_1 <= tile_7_filtered_output(23);
   bh14_w99_0 <= tile_7_filtered_output(24);
   bh14_w100_0 <= tile_7_filtered_output(25);
   bh14_w101_0 <= tile_7_filtered_output(26);
   bh14_w102_0 <= tile_7_filtered_output(27);
   bh14_w103_0 <= tile_7_filtered_output(28);
   bh14_w104_0 <= tile_7_filtered_output(29);
   bh14_w105_0 <= tile_7_filtered_output(30);
   bh14_w106_0 <= tile_7_filtered_output(31);
   bh14_w107_0 <= tile_7_filtered_output(32);
   bh14_w108_0 <= not tile_7_filtered_output(33);
   tile_8_X <= X(16 downto 0);
   tile_8_Y <= Y(60 downto 48);
   tile_8_mult: DSPBlock_17x13_F50_uid32
      port map ( clk  => clk,
                 X => tile_8_X,
                 Y => tile_8_Y,
                 R => tile_8_output);

   tile_8_filtered_output <= signed(tile_8_output(29 downto 0));
   bh14_w48_4 <= tile_8_filtered_output(0);
   bh14_w49_4 <= tile_8_filtered_output(1);
   bh14_w50_4 <= tile_8_filtered_output(2);
   bh14_w51_5 <= tile_8_filtered_output(3);
   bh14_w52_5 <= tile_8_filtered_output(4);
   bh14_w53_5 <= tile_8_filtered_output(5);
   bh14_w54_5 <= tile_8_filtered_output(6);
   bh14_w55_5 <= tile_8_filtered_output(7);
   bh14_w56_5 <= tile_8_filtered_output(8);
   bh14_w57_5 <= tile_8_filtered_output(9);
   bh14_w58_5 <= tile_8_filtered_output(10);
   bh14_w59_5 <= tile_8_filtered_output(11);
   bh14_w60_5 <= tile_8_filtered_output(12);
   bh14_w61_5 <= tile_8_filtered_output(13);
   bh14_w62_5 <= tile_8_filtered_output(14);
   bh14_w63_5 <= tile_8_filtered_output(15);
   bh14_w64_5 <= tile_8_filtered_output(16);
   bh14_w65_4 <= tile_8_filtered_output(17);
   bh14_w66_4 <= tile_8_filtered_output(18);
   bh14_w67_4 <= tile_8_filtered_output(19);
   bh14_w68_4 <= tile_8_filtered_output(20);
   bh14_w69_4 <= tile_8_filtered_output(21);
   bh14_w70_4 <= tile_8_filtered_output(22);
   bh14_w71_4 <= tile_8_filtered_output(23);
   bh14_w72_4 <= tile_8_filtered_output(24);
   bh14_w73_4 <= tile_8_filtered_output(25);
   bh14_w74_4 <= tile_8_filtered_output(26);
   bh14_w75_4 <= tile_8_filtered_output(27);
   bh14_w76_4 <= tile_8_filtered_output(28);
   bh14_w77_4 <= not tile_8_filtered_output(29);
   tile_9_X <= X(33 downto 17);
   tile_9_Y <= Y(60 downto 48);
   tile_9_mult: DSPBlock_17x13_F50_uid34
      port map ( clk  => clk,
                 X => tile_9_X,
                 Y => tile_9_Y,
                 R => tile_9_output);

   tile_9_filtered_output <= signed(tile_9_output(29 downto 0));
   bh14_w65_5 <= tile_9_filtered_output(0);
   bh14_w66_5 <= tile_9_filtered_output(1);
   bh14_w67_5 <= tile_9_filtered_output(2);
   bh14_w68_5 <= tile_9_filtered_output(3);
   bh14_w69_5 <= tile_9_filtered_output(4);
   bh14_w70_5 <= tile_9_filtered_output(5);
   bh14_w71_5 <= tile_9_filtered_output(6);
   bh14_w72_5 <= tile_9_filtered_output(7);
   bh14_w73_5 <= tile_9_filtered_output(8);
   bh14_w74_5 <= tile_9_filtered_output(9);
   bh14_w75_5 <= tile_9_filtered_output(10);
   bh14_w76_5 <= tile_9_filtered_output(11);
   bh14_w77_5 <= tile_9_filtered_output(12);
   bh14_w78_4 <= tile_9_filtered_output(13);
   bh14_w79_4 <= tile_9_filtered_output(14);
   bh14_w80_4 <= tile_9_filtered_output(15);
   bh14_w81_4 <= tile_9_filtered_output(16);
   bh14_w82_3 <= tile_9_filtered_output(17);
   bh14_w83_3 <= tile_9_filtered_output(18);
   bh14_w84_3 <= tile_9_filtered_output(19);
   bh14_w85_2 <= tile_9_filtered_output(20);
   bh14_w86_2 <= tile_9_filtered_output(21);
   bh14_w87_2 <= tile_9_filtered_output(22);
   bh14_w88_2 <= tile_9_filtered_output(23);
   bh14_w89_2 <= tile_9_filtered_output(24);
   bh14_w90_2 <= tile_9_filtered_output(25);
   bh14_w91_2 <= tile_9_filtered_output(26);
   bh14_w92_2 <= tile_9_filtered_output(27);
   bh14_w93_2 <= tile_9_filtered_output(28);
   bh14_w94_2 <= not tile_9_filtered_output(29);
   tile_10_X <= X(50 downto 34);
   tile_10_Y <= Y(60 downto 48);
   tile_10_mult: DSPBlock_17x13_F50_uid36
      port map ( clk  => clk,
                 X => tile_10_X,
                 Y => tile_10_Y,
                 R => tile_10_output);

   tile_10_filtered_output <= signed(tile_10_output(29 downto 0));
   bh14_w82_4 <= tile_10_filtered_output(0);
   bh14_w83_4 <= tile_10_filtered_output(1);
   bh14_w84_4 <= tile_10_filtered_output(2);
   bh14_w85_3 <= tile_10_filtered_output(3);
   bh14_w86_3 <= tile_10_filtered_output(4);
   bh14_w87_3 <= tile_10_filtered_output(5);
   bh14_w88_3 <= tile_10_filtered_output(6);
   bh14_w89_3 <= tile_10_filtered_output(7);
   bh14_w90_3 <= tile_10_filtered_output(8);
   bh14_w91_3 <= tile_10_filtered_output(9);
   bh14_w92_3 <= tile_10_filtered_output(10);
   bh14_w93_3 <= tile_10_filtered_output(11);
   bh14_w94_3 <= tile_10_filtered_output(12);
   bh14_w95_2 <= tile_10_filtered_output(13);
   bh14_w96_2 <= tile_10_filtered_output(14);
   bh14_w97_2 <= tile_10_filtered_output(15);
   bh14_w98_2 <= tile_10_filtered_output(16);
   bh14_w99_1 <= tile_10_filtered_output(17);
   bh14_w100_1 <= tile_10_filtered_output(18);
   bh14_w101_1 <= tile_10_filtered_output(19);
   bh14_w102_1 <= tile_10_filtered_output(20);
   bh14_w103_1 <= tile_10_filtered_output(21);
   bh14_w104_1 <= tile_10_filtered_output(22);
   bh14_w105_1 <= tile_10_filtered_output(23);
   bh14_w106_1 <= tile_10_filtered_output(24);
   bh14_w107_1 <= tile_10_filtered_output(25);
   bh14_w108_1 <= tile_10_filtered_output(26);
   bh14_w109_0 <= tile_10_filtered_output(27);
   bh14_w110_0 <= tile_10_filtered_output(28);
   bh14_w111_0 <= not tile_10_filtered_output(29);
   tile_11_X <= X(60 downto 51);
   tile_11_Y <= Y(60 downto 48);
   tile_11_mult: DSPBlock_10x13_F50_uid38
      port map ( clk  => clk,
                 X => tile_11_X,
                 Y => tile_11_Y,
                 R => tile_11_output);

   tile_11_filtered_output <= signed(tile_11_output(22 downto 0));
   bh14_w99_2 <= tile_11_filtered_output(0);
   bh14_w100_2 <= tile_11_filtered_output(1);
   bh14_w101_2 <= tile_11_filtered_output(2);
   bh14_w102_2 <= tile_11_filtered_output(3);
   bh14_w103_2 <= tile_11_filtered_output(4);
   bh14_w104_2 <= tile_11_filtered_output(5);
   bh14_w105_2 <= tile_11_filtered_output(6);
   bh14_w106_2 <= tile_11_filtered_output(7);
   bh14_w107_2 <= tile_11_filtered_output(8);
   bh14_w108_2 <= tile_11_filtered_output(9);
   bh14_w109_1 <= tile_11_filtered_output(10);
   bh14_w110_1 <= tile_11_filtered_output(11);
   bh14_w111_1 <= tile_11_filtered_output(12);
   bh14_w112_0 <= tile_11_filtered_output(13);
   bh14_w113_0 <= tile_11_filtered_output(14);
   bh14_w114_0 <= tile_11_filtered_output(15);
   bh14_w115_0 <= tile_11_filtered_output(16);
   bh14_w116_0 <= tile_11_filtered_output(17);
   bh14_w117_0 <= tile_11_filtered_output(18);
   bh14_w118_0 <= tile_11_filtered_output(19);
   bh14_w119_0 <= tile_11_filtered_output(20);
   bh14_w120_0 <= tile_11_filtered_output(21);
   bh14_w121_0 <= not tile_11_filtered_output(22);

   -- Adding the constant bits 
   bh14_w77_6 <= '1';
   bh14_w78_5 <= '1';
   bh14_w79_5 <= '1';
   bh14_w80_5 <= '1';
   bh14_w81_5 <= '1';
   bh14_w82_5 <= '1';
   bh14_w83_5 <= '1';
   bh14_w85_4 <= '1';
   bh14_w86_4 <= '1';
   bh14_w87_4 <= '1';
   bh14_w88_4 <= '1';
   bh14_w89_4 <= '1';
   bh14_w90_4 <= '1';
   bh14_w91_4 <= '1';
   bh14_w92_4 <= '1';
   bh14_w93_4 <= '1';
   bh14_w95_3 <= '1';
   bh14_w96_3 <= '1';
   bh14_w97_3 <= '1';
   bh14_w98_3 <= '1';
   bh14_w99_3 <= '1';
   bh14_w100_3 <= '1';
   bh14_w101_3 <= '1';
   bh14_w102_3 <= '1';
   bh14_w103_3 <= '1';
   bh14_w104_3 <= '1';
   bh14_w105_3 <= '1';
   bh14_w106_3 <= '1';
   bh14_w107_3 <= '1';
   bh14_w109_2 <= '1';
   bh14_w110_2 <= '1';
   bh14_w112_1 <= '1';
   bh14_w113_1 <= '1';
   bh14_w114_1 <= '1';
   bh14_w115_1 <= '1';
   bh14_w116_1 <= '1';
   bh14_w117_1 <= '1';
   bh14_w118_1 <= '1';
   bh14_w119_1 <= '1';
   bh14_w120_1 <= '1';


   Compressor_23_3_F50_uid41_bh14_uid42_In0 <= "" & bh14_w17_0 & bh14_w17_1 & "0";
   Compressor_23_3_F50_uid41_bh14_uid42_In1 <= "" & bh14_w18_0 & bh14_w18_1;
   Compressor_23_3_F50_uid41_uid42: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid42_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid42_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid42_Out0_copy43);
   Compressor_23_3_F50_uid41_bh14_uid42_Out0 <= Compressor_23_3_F50_uid41_bh14_uid42_Out0_copy43; -- output copy to hold a pipeline register if needed

   bh14_w17_2 <= Compressor_23_3_F50_uid41_bh14_uid42_Out0(0);
   bh14_w18_2 <= Compressor_23_3_F50_uid41_bh14_uid42_Out0(1);
   bh14_w19_2 <= Compressor_23_3_F50_uid41_bh14_uid42_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid44_In0 <= "" & bh14_w19_0 & bh14_w19_1 & "0";
   Compressor_23_3_F50_uid41_bh14_uid44_In1 <= "" & bh14_w20_0 & bh14_w20_1;
   Compressor_23_3_F50_uid41_uid44: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid44_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid44_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid44_Out0_copy45);
   Compressor_23_3_F50_uid41_bh14_uid44_Out0 <= Compressor_23_3_F50_uid41_bh14_uid44_Out0_copy45; -- output copy to hold a pipeline register if needed

   bh14_w19_3 <= Compressor_23_3_F50_uid41_bh14_uid44_Out0(0);
   bh14_w20_2 <= Compressor_23_3_F50_uid41_bh14_uid44_Out0(1);
   bh14_w21_2 <= Compressor_23_3_F50_uid41_bh14_uid44_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid46_In0 <= "" & bh14_w21_0 & bh14_w21_1 & "0";
   Compressor_23_3_F50_uid41_bh14_uid46_In1 <= "" & bh14_w22_0 & bh14_w22_1;
   Compressor_23_3_F50_uid41_uid46: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid46_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid46_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid46_Out0_copy47);
   Compressor_23_3_F50_uid41_bh14_uid46_Out0 <= Compressor_23_3_F50_uid41_bh14_uid46_Out0_copy47; -- output copy to hold a pipeline register if needed

   bh14_w21_3 <= Compressor_23_3_F50_uid41_bh14_uid46_Out0(0);
   bh14_w22_2 <= Compressor_23_3_F50_uid41_bh14_uid46_Out0(1);
   bh14_w23_2 <= Compressor_23_3_F50_uid41_bh14_uid46_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid50_In0 <= "" & bh14_w23_0 & bh14_w23_1 & "0";
   Compressor_3_2_F50_uid49_uid50: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid50_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid50_Out0_copy51);
   Compressor_3_2_F50_uid49_bh14_uid50_Out0 <= Compressor_3_2_F50_uid49_bh14_uid50_Out0_copy51; -- output copy to hold a pipeline register if needed

   bh14_w23_3 <= Compressor_3_2_F50_uid49_bh14_uid50_Out0(0);
   bh14_w24_3 <= Compressor_3_2_F50_uid49_bh14_uid50_Out0(1);

   Compressor_23_3_F50_uid41_bh14_uid52_In0 <= "" & bh14_w24_0 & bh14_w24_1 & bh14_w24_2;
   Compressor_23_3_F50_uid41_bh14_uid52_In1 <= "" & bh14_w25_0 & bh14_w25_1;
   Compressor_23_3_F50_uid41_uid52: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid52_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid52_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid52_Out0_copy53);
   Compressor_23_3_F50_uid41_bh14_uid52_Out0 <= Compressor_23_3_F50_uid41_bh14_uid52_Out0_copy53; -- output copy to hold a pipeline register if needed

   bh14_w24_4 <= Compressor_23_3_F50_uid41_bh14_uid52_Out0(0);
   bh14_w25_3 <= Compressor_23_3_F50_uid41_bh14_uid52_Out0(1);
   bh14_w26_3 <= Compressor_23_3_F50_uid41_bh14_uid52_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid54_In0 <= "" & bh14_w26_0 & bh14_w26_1 & bh14_w26_2;
   Compressor_23_3_F50_uid41_bh14_uid54_In1 <= "" & bh14_w27_0 & bh14_w27_1;
   Compressor_23_3_F50_uid41_uid54: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid54_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid54_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid54_Out0_copy55);
   Compressor_23_3_F50_uid41_bh14_uid54_Out0 <= Compressor_23_3_F50_uid41_bh14_uid54_Out0_copy55; -- output copy to hold a pipeline register if needed

   bh14_w26_4 <= Compressor_23_3_F50_uid41_bh14_uid54_Out0(0);
   bh14_w27_3 <= Compressor_23_3_F50_uid41_bh14_uid54_Out0(1);
   bh14_w28_3 <= Compressor_23_3_F50_uid41_bh14_uid54_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid56_In0 <= "" & bh14_w28_0 & bh14_w28_1 & bh14_w28_2;
   Compressor_23_3_F50_uid41_bh14_uid56_In1 <= "" & bh14_w29_0 & bh14_w29_1;
   Compressor_23_3_F50_uid41_uid56: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid56_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid56_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid56_Out0_copy57);
   Compressor_23_3_F50_uid41_bh14_uid56_Out0 <= Compressor_23_3_F50_uid41_bh14_uid56_Out0_copy57; -- output copy to hold a pipeline register if needed

   bh14_w28_4 <= Compressor_23_3_F50_uid41_bh14_uid56_Out0(0);
   bh14_w29_3 <= Compressor_23_3_F50_uid41_bh14_uid56_Out0(1);
   bh14_w30_3 <= Compressor_23_3_F50_uid41_bh14_uid56_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid58_In0 <= "" & bh14_w30_0 & bh14_w30_1 & bh14_w30_2;
   Compressor_23_3_F50_uid41_bh14_uid58_In1 <= "" & bh14_w31_0 & bh14_w31_1;
   Compressor_23_3_F50_uid41_uid58: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid58_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid58_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid58_Out0_copy59);
   Compressor_23_3_F50_uid41_bh14_uid58_Out0 <= Compressor_23_3_F50_uid41_bh14_uid58_Out0_copy59; -- output copy to hold a pipeline register if needed

   bh14_w30_4 <= Compressor_23_3_F50_uid41_bh14_uid58_Out0(0);
   bh14_w31_3 <= Compressor_23_3_F50_uid41_bh14_uid58_Out0(1);
   bh14_w32_3 <= Compressor_23_3_F50_uid41_bh14_uid58_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid60_In0 <= "" & bh14_w32_0 & bh14_w32_1 & bh14_w32_2;
   Compressor_23_3_F50_uid41_bh14_uid60_In1 <= "" & bh14_w33_0 & bh14_w33_1;
   Compressor_23_3_F50_uid41_uid60: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid60_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid60_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid60_Out0_copy61);
   Compressor_23_3_F50_uid41_bh14_uid60_Out0 <= Compressor_23_3_F50_uid41_bh14_uid60_Out0_copy61; -- output copy to hold a pipeline register if needed

   bh14_w32_4 <= Compressor_23_3_F50_uid41_bh14_uid60_Out0(0);
   bh14_w33_3 <= Compressor_23_3_F50_uid41_bh14_uid60_Out0(1);
   bh14_w34_4 <= Compressor_23_3_F50_uid41_bh14_uid60_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid64_In0 <= "" & bh14_w34_0 & bh14_w34_1 & bh14_w34_2 & bh14_w34_3;
   Compressor_14_3_F50_uid63_bh14_uid64_In1 <= "" & bh14_w35_0;
   Compressor_14_3_F50_uid63_uid64: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid64_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid64_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid64_Out0_copy65);
   Compressor_14_3_F50_uid63_bh14_uid64_Out0 <= Compressor_14_3_F50_uid63_bh14_uid64_Out0_copy65; -- output copy to hold a pipeline register if needed

   bh14_w34_5 <= Compressor_14_3_F50_uid63_bh14_uid64_Out0(0);
   bh14_w35_4 <= Compressor_14_3_F50_uid63_bh14_uid64_Out0(1);
   bh14_w36_4 <= Compressor_14_3_F50_uid63_bh14_uid64_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid66_In0 <= "" & bh14_w35_1 & bh14_w35_2 & bh14_w35_3;
   Compressor_3_2_F50_uid49_uid66: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid66_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid66_Out0_copy67);
   Compressor_3_2_F50_uid49_bh14_uid66_Out0 <= Compressor_3_2_F50_uid49_bh14_uid66_Out0_copy67; -- output copy to hold a pipeline register if needed

   bh14_w35_5 <= Compressor_3_2_F50_uid49_bh14_uid66_Out0(0);
   bh14_w36_5 <= Compressor_3_2_F50_uid49_bh14_uid66_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid68_In0 <= "" & bh14_w36_0 & bh14_w36_1 & bh14_w36_2 & bh14_w36_3;
   Compressor_14_3_F50_uid63_bh14_uid68_In1 <= "" & bh14_w37_0;
   Compressor_14_3_F50_uid63_uid68: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid68_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid68_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid68_Out0_copy69);
   Compressor_14_3_F50_uid63_bh14_uid68_Out0 <= Compressor_14_3_F50_uid63_bh14_uid68_Out0_copy69; -- output copy to hold a pipeline register if needed

   bh14_w36_6 <= Compressor_14_3_F50_uid63_bh14_uid68_Out0(0);
   bh14_w37_4 <= Compressor_14_3_F50_uid63_bh14_uid68_Out0(1);
   bh14_w38_4 <= Compressor_14_3_F50_uid63_bh14_uid68_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid70_In0 <= "" & bh14_w37_1 & bh14_w37_2 & bh14_w37_3;
   Compressor_3_2_F50_uid49_uid70: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid70_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid70_Out0_copy71);
   Compressor_3_2_F50_uid49_bh14_uid70_Out0 <= Compressor_3_2_F50_uid49_bh14_uid70_Out0_copy71; -- output copy to hold a pipeline register if needed

   bh14_w37_5 <= Compressor_3_2_F50_uid49_bh14_uid70_Out0(0);
   bh14_w38_5 <= Compressor_3_2_F50_uid49_bh14_uid70_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid72_In0 <= "" & bh14_w38_0 & bh14_w38_1 & bh14_w38_2 & bh14_w38_3;
   Compressor_14_3_F50_uid63_bh14_uid72_In1 <= "" & bh14_w39_0;
   Compressor_14_3_F50_uid63_uid72: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid72_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid72_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid72_Out0_copy73);
   Compressor_14_3_F50_uid63_bh14_uid72_Out0 <= Compressor_14_3_F50_uid63_bh14_uid72_Out0_copy73; -- output copy to hold a pipeline register if needed

   bh14_w38_6 <= Compressor_14_3_F50_uid63_bh14_uid72_Out0(0);
   bh14_w39_4 <= Compressor_14_3_F50_uid63_bh14_uid72_Out0(1);
   bh14_w40_4 <= Compressor_14_3_F50_uid63_bh14_uid72_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid74_In0 <= "" & bh14_w39_1 & bh14_w39_2 & bh14_w39_3;
   Compressor_3_2_F50_uid49_uid74: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid74_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid74_Out0_copy75);
   Compressor_3_2_F50_uid49_bh14_uid74_Out0 <= Compressor_3_2_F50_uid49_bh14_uid74_Out0_copy75; -- output copy to hold a pipeline register if needed

   bh14_w39_5 <= Compressor_3_2_F50_uid49_bh14_uid74_Out0(0);
   bh14_w40_5 <= Compressor_3_2_F50_uid49_bh14_uid74_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid76_In0 <= "" & bh14_w40_0 & bh14_w40_1 & bh14_w40_2 & bh14_w40_3;
   Compressor_14_3_F50_uid63_bh14_uid76_In1 <= "" & bh14_w41_0;
   Compressor_14_3_F50_uid63_uid76: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid76_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid76_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid76_Out0_copy77);
   Compressor_14_3_F50_uid63_bh14_uid76_Out0 <= Compressor_14_3_F50_uid63_bh14_uid76_Out0_copy77; -- output copy to hold a pipeline register if needed

   bh14_w40_6 <= Compressor_14_3_F50_uid63_bh14_uid76_Out0(0);
   bh14_w41_4 <= Compressor_14_3_F50_uid63_bh14_uid76_Out0(1);
   bh14_w42_4 <= Compressor_14_3_F50_uid63_bh14_uid76_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid78_In0 <= "" & bh14_w41_1 & bh14_w41_2 & bh14_w41_3;
   Compressor_3_2_F50_uid49_uid78: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid78_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid78_Out0_copy79);
   Compressor_3_2_F50_uid49_bh14_uid78_Out0 <= Compressor_3_2_F50_uid49_bh14_uid78_Out0_copy79; -- output copy to hold a pipeline register if needed

   bh14_w41_5 <= Compressor_3_2_F50_uid49_bh14_uid78_Out0(0);
   bh14_w42_5 <= Compressor_3_2_F50_uid49_bh14_uid78_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid80_In0 <= "" & bh14_w42_0 & bh14_w42_1 & bh14_w42_2 & bh14_w42_3;
   Compressor_14_3_F50_uid63_bh14_uid80_In1 <= "" & bh14_w43_0;
   Compressor_14_3_F50_uid63_uid80: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid80_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid80_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid80_Out0_copy81);
   Compressor_14_3_F50_uid63_bh14_uid80_Out0 <= Compressor_14_3_F50_uid63_bh14_uid80_Out0_copy81; -- output copy to hold a pipeline register if needed

   bh14_w42_6 <= Compressor_14_3_F50_uid63_bh14_uid80_Out0(0);
   bh14_w43_4 <= Compressor_14_3_F50_uid63_bh14_uid80_Out0(1);
   bh14_w44_4 <= Compressor_14_3_F50_uid63_bh14_uid80_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid82_In0 <= "" & bh14_w43_1 & bh14_w43_2 & bh14_w43_3;
   Compressor_3_2_F50_uid49_uid82: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid82_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid82_Out0_copy83);
   Compressor_3_2_F50_uid49_bh14_uid82_Out0 <= Compressor_3_2_F50_uid49_bh14_uid82_Out0_copy83; -- output copy to hold a pipeline register if needed

   bh14_w43_5 <= Compressor_3_2_F50_uid49_bh14_uid82_Out0(0);
   bh14_w44_5 <= Compressor_3_2_F50_uid49_bh14_uid82_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid84_In0 <= "" & bh14_w44_0 & bh14_w44_1 & bh14_w44_2 & bh14_w44_3;
   Compressor_14_3_F50_uid63_bh14_uid84_In1 <= "" & bh14_w45_0;
   Compressor_14_3_F50_uid63_uid84: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid84_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid84_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid84_Out0_copy85);
   Compressor_14_3_F50_uid63_bh14_uid84_Out0 <= Compressor_14_3_F50_uid63_bh14_uid84_Out0_copy85; -- output copy to hold a pipeline register if needed

   bh14_w44_6 <= Compressor_14_3_F50_uid63_bh14_uid84_Out0(0);
   bh14_w45_4 <= Compressor_14_3_F50_uid63_bh14_uid84_Out0(1);
   bh14_w46_4 <= Compressor_14_3_F50_uid63_bh14_uid84_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid86_In0 <= "" & bh14_w45_1 & bh14_w45_2 & bh14_w45_3;
   Compressor_3_2_F50_uid49_uid86: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid86_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid86_Out0_copy87);
   Compressor_3_2_F50_uid49_bh14_uid86_Out0 <= Compressor_3_2_F50_uid49_bh14_uid86_Out0_copy87; -- output copy to hold a pipeline register if needed

   bh14_w45_5 <= Compressor_3_2_F50_uid49_bh14_uid86_Out0(0);
   bh14_w46_5 <= Compressor_3_2_F50_uid49_bh14_uid86_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid88_In0 <= "" & bh14_w46_0 & bh14_w46_1 & bh14_w46_2 & bh14_w46_3;
   Compressor_14_3_F50_uid63_bh14_uid88_In1 <= "" & bh14_w47_0;
   Compressor_14_3_F50_uid63_uid88: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid88_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid88_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid88_Out0_copy89);
   Compressor_14_3_F50_uid63_bh14_uid88_Out0 <= Compressor_14_3_F50_uid63_bh14_uid88_Out0_copy89; -- output copy to hold a pipeline register if needed

   bh14_w46_6 <= Compressor_14_3_F50_uid63_bh14_uid88_Out0(0);
   bh14_w47_4 <= Compressor_14_3_F50_uid63_bh14_uid88_Out0(1);
   bh14_w48_5 <= Compressor_14_3_F50_uid63_bh14_uid88_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid90_In0 <= "" & bh14_w47_1 & bh14_w47_2 & bh14_w47_3;
   Compressor_3_2_F50_uid49_uid90: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid90_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid90_Out0_copy91);
   Compressor_3_2_F50_uid49_bh14_uid90_Out0 <= Compressor_3_2_F50_uid49_bh14_uid90_Out0_copy91; -- output copy to hold a pipeline register if needed

   bh14_w47_5 <= Compressor_3_2_F50_uid49_bh14_uid90_Out0(0);
   bh14_w48_6 <= Compressor_3_2_F50_uid49_bh14_uid90_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid92_In0 <= "" & bh14_w48_0 & bh14_w48_1 & bh14_w48_2 & bh14_w48_3;
   Compressor_14_3_F50_uid63_bh14_uid92_In1 <= "" & bh14_w49_0;
   Compressor_14_3_F50_uid63_uid92: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid92_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid92_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid92_Out0_copy93);
   Compressor_14_3_F50_uid63_bh14_uid92_Out0 <= Compressor_14_3_F50_uid63_bh14_uid92_Out0_copy93; -- output copy to hold a pipeline register if needed

   bh14_w48_7 <= Compressor_14_3_F50_uid63_bh14_uid92_Out0(0);
   bh14_w49_5 <= Compressor_14_3_F50_uid63_bh14_uid92_Out0(1);
   bh14_w50_5 <= Compressor_14_3_F50_uid63_bh14_uid92_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid94_In0 <= "" & bh14_w49_1 & bh14_w49_2 & bh14_w49_3 & bh14_w49_4;
   Compressor_14_3_F50_uid63_bh14_uid94_In1 <= "" & bh14_w50_0;
   Compressor_14_3_F50_uid63_uid94: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid94_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid94_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid94_Out0_copy95);
   Compressor_14_3_F50_uid63_bh14_uid94_Out0 <= Compressor_14_3_F50_uid63_bh14_uid94_Out0_copy95; -- output copy to hold a pipeline register if needed

   bh14_w49_6 <= Compressor_14_3_F50_uid63_bh14_uid94_Out0(0);
   bh14_w50_6 <= Compressor_14_3_F50_uid63_bh14_uid94_Out0(1);
   bh14_w51_6 <= Compressor_14_3_F50_uid63_bh14_uid94_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid96_In0 <= "" & bh14_w50_1 & bh14_w50_2 & bh14_w50_3;
   Compressor_3_2_F50_uid49_uid96: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid96_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid96_Out0_copy97);
   Compressor_3_2_F50_uid49_bh14_uid96_Out0 <= Compressor_3_2_F50_uid49_bh14_uid96_Out0_copy97; -- output copy to hold a pipeline register if needed

   bh14_w50_7 <= Compressor_3_2_F50_uid49_bh14_uid96_Out0(0);
   bh14_w51_7 <= Compressor_3_2_F50_uid49_bh14_uid96_Out0(1);

   Compressor_6_3_F50_uid99_bh14_uid100_In0 <= "" & bh14_w51_0 & bh14_w51_1 & bh14_w51_2 & bh14_w51_3 & bh14_w51_4 & bh14_w51_5;
   Compressor_6_3_F50_uid99_uid100: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid100_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid100_Out0_copy101);
   Compressor_6_3_F50_uid99_bh14_uid100_Out0 <= Compressor_6_3_F50_uid99_bh14_uid100_Out0_copy101; -- output copy to hold a pipeline register if needed

   bh14_w51_8 <= Compressor_6_3_F50_uid99_bh14_uid100_Out0(0);
   bh14_w52_6 <= Compressor_6_3_F50_uid99_bh14_uid100_Out0(1);
   bh14_w53_6 <= Compressor_6_3_F50_uid99_bh14_uid100_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid102_In0 <= "" & bh14_w52_0 & bh14_w52_1 & bh14_w52_2 & bh14_w52_3 & bh14_w52_4 & bh14_w52_5;
   Compressor_6_3_F50_uid99_uid102: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid102_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid102_Out0_copy103);
   Compressor_6_3_F50_uid99_bh14_uid102_Out0 <= Compressor_6_3_F50_uid99_bh14_uid102_Out0_copy103; -- output copy to hold a pipeline register if needed

   bh14_w52_7 <= Compressor_6_3_F50_uid99_bh14_uid102_Out0(0);
   bh14_w53_7 <= Compressor_6_3_F50_uid99_bh14_uid102_Out0(1);
   bh14_w54_6 <= Compressor_6_3_F50_uid99_bh14_uid102_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid104_In0 <= "" & bh14_w53_0 & bh14_w53_1 & bh14_w53_2 & bh14_w53_3 & bh14_w53_4 & bh14_w53_5;
   Compressor_6_3_F50_uid99_uid104: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid104_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid104_Out0_copy105);
   Compressor_6_3_F50_uid99_bh14_uid104_Out0 <= Compressor_6_3_F50_uid99_bh14_uid104_Out0_copy105; -- output copy to hold a pipeline register if needed

   bh14_w53_8 <= Compressor_6_3_F50_uid99_bh14_uid104_Out0(0);
   bh14_w54_7 <= Compressor_6_3_F50_uid99_bh14_uid104_Out0(1);
   bh14_w55_6 <= Compressor_6_3_F50_uid99_bh14_uid104_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid106_In0 <= "" & bh14_w54_0 & bh14_w54_1 & bh14_w54_2 & bh14_w54_3 & bh14_w54_4 & bh14_w54_5;
   Compressor_6_3_F50_uid99_uid106: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid106_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid106_Out0_copy107);
   Compressor_6_3_F50_uid99_bh14_uid106_Out0 <= Compressor_6_3_F50_uid99_bh14_uid106_Out0_copy107; -- output copy to hold a pipeline register if needed

   bh14_w54_8 <= Compressor_6_3_F50_uid99_bh14_uid106_Out0(0);
   bh14_w55_7 <= Compressor_6_3_F50_uid99_bh14_uid106_Out0(1);
   bh14_w56_6 <= Compressor_6_3_F50_uid99_bh14_uid106_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid108_In0 <= "" & bh14_w55_0 & bh14_w55_1 & bh14_w55_2 & bh14_w55_3 & bh14_w55_4 & bh14_w55_5;
   Compressor_6_3_F50_uid99_uid108: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid108_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid108_Out0_copy109);
   Compressor_6_3_F50_uid99_bh14_uid108_Out0 <= Compressor_6_3_F50_uid99_bh14_uid108_Out0_copy109; -- output copy to hold a pipeline register if needed

   bh14_w55_8 <= Compressor_6_3_F50_uid99_bh14_uid108_Out0(0);
   bh14_w56_7 <= Compressor_6_3_F50_uid99_bh14_uid108_Out0(1);
   bh14_w57_6 <= Compressor_6_3_F50_uid99_bh14_uid108_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid110_In0 <= "" & bh14_w56_0 & bh14_w56_1 & bh14_w56_2 & bh14_w56_3 & bh14_w56_4 & bh14_w56_5;
   Compressor_6_3_F50_uid99_uid110: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid110_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid110_Out0_copy111);
   Compressor_6_3_F50_uid99_bh14_uid110_Out0 <= Compressor_6_3_F50_uid99_bh14_uid110_Out0_copy111; -- output copy to hold a pipeline register if needed

   bh14_w56_8 <= Compressor_6_3_F50_uid99_bh14_uid110_Out0(0);
   bh14_w57_7 <= Compressor_6_3_F50_uid99_bh14_uid110_Out0(1);
   bh14_w58_6 <= Compressor_6_3_F50_uid99_bh14_uid110_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid112_In0 <= "" & bh14_w57_0 & bh14_w57_1 & bh14_w57_2 & bh14_w57_3 & bh14_w57_4 & bh14_w57_5;
   Compressor_6_3_F50_uid99_uid112: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid112_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid112_Out0_copy113);
   Compressor_6_3_F50_uid99_bh14_uid112_Out0 <= Compressor_6_3_F50_uid99_bh14_uid112_Out0_copy113; -- output copy to hold a pipeline register if needed

   bh14_w57_8 <= Compressor_6_3_F50_uid99_bh14_uid112_Out0(0);
   bh14_w58_7 <= Compressor_6_3_F50_uid99_bh14_uid112_Out0(1);
   bh14_w59_6 <= Compressor_6_3_F50_uid99_bh14_uid112_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid114_In0 <= "" & bh14_w58_0 & bh14_w58_1 & bh14_w58_2 & bh14_w58_3 & bh14_w58_4 & bh14_w58_5;
   Compressor_6_3_F50_uid99_uid114: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid114_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid114_Out0_copy115);
   Compressor_6_3_F50_uid99_bh14_uid114_Out0 <= Compressor_6_3_F50_uid99_bh14_uid114_Out0_copy115; -- output copy to hold a pipeline register if needed

   bh14_w58_8 <= Compressor_6_3_F50_uid99_bh14_uid114_Out0(0);
   bh14_w59_7 <= Compressor_6_3_F50_uid99_bh14_uid114_Out0(1);
   bh14_w60_6 <= Compressor_6_3_F50_uid99_bh14_uid114_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid116_In0 <= "" & bh14_w59_0 & bh14_w59_1 & bh14_w59_2 & bh14_w59_3 & bh14_w59_4 & bh14_w59_5;
   Compressor_6_3_F50_uid99_uid116: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid116_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid116_Out0_copy117);
   Compressor_6_3_F50_uid99_bh14_uid116_Out0 <= Compressor_6_3_F50_uid99_bh14_uid116_Out0_copy117; -- output copy to hold a pipeline register if needed

   bh14_w59_8 <= Compressor_6_3_F50_uid99_bh14_uid116_Out0(0);
   bh14_w60_7 <= Compressor_6_3_F50_uid99_bh14_uid116_Out0(1);
   bh14_w61_6 <= Compressor_6_3_F50_uid99_bh14_uid116_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid118_In0 <= "" & bh14_w60_0 & bh14_w60_1 & bh14_w60_2 & bh14_w60_3 & bh14_w60_4 & bh14_w60_5;
   Compressor_6_3_F50_uid99_uid118: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid118_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid118_Out0_copy119);
   Compressor_6_3_F50_uid99_bh14_uid118_Out0 <= Compressor_6_3_F50_uid99_bh14_uid118_Out0_copy119; -- output copy to hold a pipeline register if needed

   bh14_w60_8 <= Compressor_6_3_F50_uid99_bh14_uid118_Out0(0);
   bh14_w61_7 <= Compressor_6_3_F50_uid99_bh14_uid118_Out0(1);
   bh14_w62_6 <= Compressor_6_3_F50_uid99_bh14_uid118_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid120_In0 <= "" & bh14_w61_0 & bh14_w61_1 & bh14_w61_2 & bh14_w61_3 & bh14_w61_4 & bh14_w61_5;
   Compressor_6_3_F50_uid99_uid120: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid120_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid120_Out0_copy121);
   Compressor_6_3_F50_uid99_bh14_uid120_Out0 <= Compressor_6_3_F50_uid99_bh14_uid120_Out0_copy121; -- output copy to hold a pipeline register if needed

   bh14_w61_8 <= Compressor_6_3_F50_uid99_bh14_uid120_Out0(0);
   bh14_w62_7 <= Compressor_6_3_F50_uid99_bh14_uid120_Out0(1);
   bh14_w63_6 <= Compressor_6_3_F50_uid99_bh14_uid120_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid122_In0 <= "" & bh14_w62_0 & bh14_w62_1 & bh14_w62_2 & bh14_w62_3 & bh14_w62_4 & bh14_w62_5;
   Compressor_6_3_F50_uid99_uid122: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid122_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid122_Out0_copy123);
   Compressor_6_3_F50_uid99_bh14_uid122_Out0 <= Compressor_6_3_F50_uid99_bh14_uid122_Out0_copy123; -- output copy to hold a pipeline register if needed

   bh14_w62_8 <= Compressor_6_3_F50_uid99_bh14_uid122_Out0(0);
   bh14_w63_7 <= Compressor_6_3_F50_uid99_bh14_uid122_Out0(1);
   bh14_w64_6 <= Compressor_6_3_F50_uid99_bh14_uid122_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid124_In0 <= "" & bh14_w63_0 & bh14_w63_1 & bh14_w63_2 & bh14_w63_3 & bh14_w63_4 & bh14_w63_5;
   Compressor_6_3_F50_uid99_uid124: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid124_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid124_Out0_copy125);
   Compressor_6_3_F50_uid99_bh14_uid124_Out0 <= Compressor_6_3_F50_uid99_bh14_uid124_Out0_copy125; -- output copy to hold a pipeline register if needed

   bh14_w63_8 <= Compressor_6_3_F50_uid99_bh14_uid124_Out0(0);
   bh14_w64_7 <= Compressor_6_3_F50_uid99_bh14_uid124_Out0(1);
   bh14_w65_6 <= Compressor_6_3_F50_uid99_bh14_uid124_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid126_In0 <= "" & bh14_w64_0 & bh14_w64_1 & bh14_w64_2 & bh14_w64_3 & bh14_w64_4 & bh14_w64_5;
   Compressor_6_3_F50_uid99_uid126: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid126_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid126_Out0_copy127);
   Compressor_6_3_F50_uid99_bh14_uid126_Out0 <= Compressor_6_3_F50_uid99_bh14_uid126_Out0_copy127; -- output copy to hold a pipeline register if needed

   bh14_w64_8 <= Compressor_6_3_F50_uid99_bh14_uid126_Out0(0);
   bh14_w65_7 <= Compressor_6_3_F50_uid99_bh14_uid126_Out0(1);
   bh14_w66_6 <= Compressor_6_3_F50_uid99_bh14_uid126_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid128_In0 <= "" & bh14_w65_0 & bh14_w65_1 & bh14_w65_2 & bh14_w65_3 & bh14_w65_4 & bh14_w65_5;
   Compressor_6_3_F50_uid99_uid128: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid128_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid128_Out0_copy129);
   Compressor_6_3_F50_uid99_bh14_uid128_Out0 <= Compressor_6_3_F50_uid99_bh14_uid128_Out0_copy129; -- output copy to hold a pipeline register if needed

   bh14_w65_8 <= Compressor_6_3_F50_uid99_bh14_uid128_Out0(0);
   bh14_w66_7 <= Compressor_6_3_F50_uid99_bh14_uid128_Out0(1);
   bh14_w67_6 <= Compressor_6_3_F50_uid99_bh14_uid128_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid130_In0 <= "" & bh14_w66_0 & bh14_w66_1 & bh14_w66_2 & bh14_w66_3 & bh14_w66_4 & bh14_w66_5;
   Compressor_6_3_F50_uid99_uid130: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid130_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid130_Out0_copy131);
   Compressor_6_3_F50_uid99_bh14_uid130_Out0 <= Compressor_6_3_F50_uid99_bh14_uid130_Out0_copy131; -- output copy to hold a pipeline register if needed

   bh14_w66_8 <= Compressor_6_3_F50_uid99_bh14_uid130_Out0(0);
   bh14_w67_7 <= Compressor_6_3_F50_uid99_bh14_uid130_Out0(1);
   bh14_w68_6 <= Compressor_6_3_F50_uid99_bh14_uid130_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid132_In0 <= "" & bh14_w67_0 & bh14_w67_1 & bh14_w67_2 & bh14_w67_3 & bh14_w67_4 & bh14_w67_5;
   Compressor_6_3_F50_uid99_uid132: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid132_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid132_Out0_copy133);
   Compressor_6_3_F50_uid99_bh14_uid132_Out0 <= Compressor_6_3_F50_uid99_bh14_uid132_Out0_copy133; -- output copy to hold a pipeline register if needed

   bh14_w67_8 <= Compressor_6_3_F50_uid99_bh14_uid132_Out0(0);
   bh14_w68_7 <= Compressor_6_3_F50_uid99_bh14_uid132_Out0(1);
   bh14_w69_6 <= Compressor_6_3_F50_uid99_bh14_uid132_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid134_In0 <= "" & bh14_w68_0 & bh14_w68_1 & bh14_w68_2 & bh14_w68_3 & bh14_w68_4 & bh14_w68_5;
   Compressor_6_3_F50_uid99_uid134: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid134_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid134_Out0_copy135);
   Compressor_6_3_F50_uid99_bh14_uid134_Out0 <= Compressor_6_3_F50_uid99_bh14_uid134_Out0_copy135; -- output copy to hold a pipeline register if needed

   bh14_w68_8 <= Compressor_6_3_F50_uid99_bh14_uid134_Out0(0);
   bh14_w69_7 <= Compressor_6_3_F50_uid99_bh14_uid134_Out0(1);
   bh14_w70_6 <= Compressor_6_3_F50_uid99_bh14_uid134_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid136_In0 <= "" & bh14_w69_0 & bh14_w69_1 & bh14_w69_2 & bh14_w69_3 & bh14_w69_4 & bh14_w69_5;
   Compressor_6_3_F50_uid99_uid136: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid136_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid136_Out0_copy137);
   Compressor_6_3_F50_uid99_bh14_uid136_Out0 <= Compressor_6_3_F50_uid99_bh14_uid136_Out0_copy137; -- output copy to hold a pipeline register if needed

   bh14_w69_8 <= Compressor_6_3_F50_uid99_bh14_uid136_Out0(0);
   bh14_w70_7 <= Compressor_6_3_F50_uid99_bh14_uid136_Out0(1);
   bh14_w71_6 <= Compressor_6_3_F50_uid99_bh14_uid136_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid138_In0 <= "" & bh14_w70_0 & bh14_w70_1 & bh14_w70_2 & bh14_w70_3 & bh14_w70_4 & bh14_w70_5;
   Compressor_6_3_F50_uid99_uid138: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid138_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid138_Out0_copy139);
   Compressor_6_3_F50_uid99_bh14_uid138_Out0 <= Compressor_6_3_F50_uid99_bh14_uid138_Out0_copy139; -- output copy to hold a pipeline register if needed

   bh14_w70_8 <= Compressor_6_3_F50_uid99_bh14_uid138_Out0(0);
   bh14_w71_7 <= Compressor_6_3_F50_uid99_bh14_uid138_Out0(1);
   bh14_w72_6 <= Compressor_6_3_F50_uid99_bh14_uid138_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid140_In0 <= "" & bh14_w71_0 & bh14_w71_1 & bh14_w71_2 & bh14_w71_3 & bh14_w71_4 & bh14_w71_5;
   Compressor_6_3_F50_uid99_uid140: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid140_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid140_Out0_copy141);
   Compressor_6_3_F50_uid99_bh14_uid140_Out0 <= Compressor_6_3_F50_uid99_bh14_uid140_Out0_copy141; -- output copy to hold a pipeline register if needed

   bh14_w71_8 <= Compressor_6_3_F50_uid99_bh14_uid140_Out0(0);
   bh14_w72_7 <= Compressor_6_3_F50_uid99_bh14_uid140_Out0(1);
   bh14_w73_6 <= Compressor_6_3_F50_uid99_bh14_uid140_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid142_In0 <= "" & bh14_w72_0 & bh14_w72_1 & bh14_w72_2 & bh14_w72_3 & bh14_w72_4 & bh14_w72_5;
   Compressor_6_3_F50_uid99_uid142: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid142_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid142_Out0_copy143);
   Compressor_6_3_F50_uid99_bh14_uid142_Out0 <= Compressor_6_3_F50_uid99_bh14_uid142_Out0_copy143; -- output copy to hold a pipeline register if needed

   bh14_w72_8 <= Compressor_6_3_F50_uid99_bh14_uid142_Out0(0);
   bh14_w73_7 <= Compressor_6_3_F50_uid99_bh14_uid142_Out0(1);
   bh14_w74_6 <= Compressor_6_3_F50_uid99_bh14_uid142_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid144_In0 <= "" & bh14_w73_0 & bh14_w73_1 & bh14_w73_2 & bh14_w73_3 & bh14_w73_4 & bh14_w73_5;
   Compressor_6_3_F50_uid99_uid144: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid144_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid144_Out0_copy145);
   Compressor_6_3_F50_uid99_bh14_uid144_Out0 <= Compressor_6_3_F50_uid99_bh14_uid144_Out0_copy145; -- output copy to hold a pipeline register if needed

   bh14_w73_8 <= Compressor_6_3_F50_uid99_bh14_uid144_Out0(0);
   bh14_w74_7 <= Compressor_6_3_F50_uid99_bh14_uid144_Out0(1);
   bh14_w75_6 <= Compressor_6_3_F50_uid99_bh14_uid144_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid146_In0 <= "" & bh14_w74_0 & bh14_w74_1 & bh14_w74_2 & bh14_w74_3 & bh14_w74_4 & bh14_w74_5;
   Compressor_6_3_F50_uid99_uid146: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid146_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid146_Out0_copy147);
   Compressor_6_3_F50_uid99_bh14_uid146_Out0 <= Compressor_6_3_F50_uid99_bh14_uid146_Out0_copy147; -- output copy to hold a pipeline register if needed

   bh14_w74_8 <= Compressor_6_3_F50_uid99_bh14_uid146_Out0(0);
   bh14_w75_7 <= Compressor_6_3_F50_uid99_bh14_uid146_Out0(1);
   bh14_w76_6 <= Compressor_6_3_F50_uid99_bh14_uid146_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid148_In0 <= "" & bh14_w75_0 & bh14_w75_1 & bh14_w75_2 & bh14_w75_3 & bh14_w75_4 & bh14_w75_5;
   Compressor_6_3_F50_uid99_uid148: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid148_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid148_Out0_copy149);
   Compressor_6_3_F50_uid99_bh14_uid148_Out0 <= Compressor_6_3_F50_uid99_bh14_uid148_Out0_copy149; -- output copy to hold a pipeline register if needed

   bh14_w75_8 <= Compressor_6_3_F50_uid99_bh14_uid148_Out0(0);
   bh14_w76_7 <= Compressor_6_3_F50_uid99_bh14_uid148_Out0(1);
   bh14_w77_7 <= Compressor_6_3_F50_uid99_bh14_uid148_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid150_In0 <= "" & bh14_w76_0 & bh14_w76_1 & bh14_w76_2 & bh14_w76_3 & bh14_w76_4 & bh14_w76_5;
   Compressor_6_3_F50_uid99_uid150: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid150_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid150_Out0_copy151);
   Compressor_6_3_F50_uid99_bh14_uid150_Out0 <= Compressor_6_3_F50_uid99_bh14_uid150_Out0_copy151; -- output copy to hold a pipeline register if needed

   bh14_w76_8 <= Compressor_6_3_F50_uid99_bh14_uid150_Out0(0);
   bh14_w77_8 <= Compressor_6_3_F50_uid99_bh14_uid150_Out0(1);
   bh14_w78_6 <= Compressor_6_3_F50_uid99_bh14_uid150_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid152_In0 <= "" & bh14_w77_0 & bh14_w77_1 & bh14_w77_2 & bh14_w77_3 & bh14_w77_4 & bh14_w77_5;
   Compressor_6_3_F50_uid99_uid152: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid152_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid152_Out0_copy153);
   Compressor_6_3_F50_uid99_bh14_uid152_Out0 <= Compressor_6_3_F50_uid99_bh14_uid152_Out0_copy153; -- output copy to hold a pipeline register if needed

   bh14_w77_9 <= Compressor_6_3_F50_uid99_bh14_uid152_Out0(0);
   bh14_w78_7 <= Compressor_6_3_F50_uid99_bh14_uid152_Out0(1);
   bh14_w79_6 <= Compressor_6_3_F50_uid99_bh14_uid152_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid154_In0 <= "" & bh14_w78_0 & bh14_w78_1 & bh14_w78_2 & bh14_w78_3 & bh14_w78_4 & bh14_w78_5;
   Compressor_6_3_F50_uid99_uid154: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid154_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid154_Out0_copy155);
   Compressor_6_3_F50_uid99_bh14_uid154_Out0 <= Compressor_6_3_F50_uid99_bh14_uid154_Out0_copy155; -- output copy to hold a pipeline register if needed

   bh14_w78_8 <= Compressor_6_3_F50_uid99_bh14_uid154_Out0(0);
   bh14_w79_7 <= Compressor_6_3_F50_uid99_bh14_uid154_Out0(1);
   bh14_w80_6 <= Compressor_6_3_F50_uid99_bh14_uid154_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid156_In0 <= "" & bh14_w79_0 & bh14_w79_1 & bh14_w79_2 & bh14_w79_3 & bh14_w79_4 & bh14_w79_5;
   Compressor_6_3_F50_uid99_uid156: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid156_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid156_Out0_copy157);
   Compressor_6_3_F50_uid99_bh14_uid156_Out0 <= Compressor_6_3_F50_uid99_bh14_uid156_Out0_copy157; -- output copy to hold a pipeline register if needed

   bh14_w79_8 <= Compressor_6_3_F50_uid99_bh14_uid156_Out0(0);
   bh14_w80_7 <= Compressor_6_3_F50_uid99_bh14_uid156_Out0(1);
   bh14_w81_6 <= Compressor_6_3_F50_uid99_bh14_uid156_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid158_In0 <= "" & bh14_w80_0 & bh14_w80_1 & bh14_w80_2 & bh14_w80_3 & bh14_w80_4 & bh14_w80_5;
   Compressor_6_3_F50_uid99_uid158: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid158_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid158_Out0_copy159);
   Compressor_6_3_F50_uid99_bh14_uid158_Out0 <= Compressor_6_3_F50_uid99_bh14_uid158_Out0_copy159; -- output copy to hold a pipeline register if needed

   bh14_w80_8 <= Compressor_6_3_F50_uid99_bh14_uid158_Out0(0);
   bh14_w81_7 <= Compressor_6_3_F50_uid99_bh14_uid158_Out0(1);
   bh14_w82_6 <= Compressor_6_3_F50_uid99_bh14_uid158_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid160_In0 <= "" & bh14_w81_0 & bh14_w81_1 & bh14_w81_2 & bh14_w81_3 & bh14_w81_4 & bh14_w81_5;
   Compressor_6_3_F50_uid99_uid160: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid160_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid160_Out0_copy161);
   Compressor_6_3_F50_uid99_bh14_uid160_Out0 <= Compressor_6_3_F50_uid99_bh14_uid160_Out0_copy161; -- output copy to hold a pipeline register if needed

   bh14_w81_8 <= Compressor_6_3_F50_uid99_bh14_uid160_Out0(0);
   bh14_w82_7 <= Compressor_6_3_F50_uid99_bh14_uid160_Out0(1);
   bh14_w83_6 <= Compressor_6_3_F50_uid99_bh14_uid160_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid162_In0 <= "" & bh14_w82_0 & bh14_w82_1 & bh14_w82_2 & bh14_w82_3 & bh14_w82_4 & bh14_w82_5;
   Compressor_6_3_F50_uid99_uid162: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid162_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid162_Out0_copy163);
   Compressor_6_3_F50_uid99_bh14_uid162_Out0 <= Compressor_6_3_F50_uid99_bh14_uid162_Out0_copy163; -- output copy to hold a pipeline register if needed

   bh14_w82_8 <= Compressor_6_3_F50_uid99_bh14_uid162_Out0(0);
   bh14_w83_7 <= Compressor_6_3_F50_uid99_bh14_uid162_Out0(1);
   bh14_w84_5 <= Compressor_6_3_F50_uid99_bh14_uid162_Out0(2);

   Compressor_6_3_F50_uid99_bh14_uid164_In0 <= "" & bh14_w83_0 & bh14_w83_1 & bh14_w83_2 & bh14_w83_3 & bh14_w83_4 & bh14_w83_5;
   Compressor_6_3_F50_uid99_uid164: Compressor_6_3_F50_uid99
      port map ( X0 => Compressor_6_3_F50_uid99_bh14_uid164_In0,
                 R => Compressor_6_3_F50_uid99_bh14_uid164_Out0_copy165);
   Compressor_6_3_F50_uid99_bh14_uid164_Out0 <= Compressor_6_3_F50_uid99_bh14_uid164_Out0_copy165; -- output copy to hold a pipeline register if needed

   bh14_w83_8 <= Compressor_6_3_F50_uid99_bh14_uid164_Out0(0);
   bh14_w84_6 <= Compressor_6_3_F50_uid99_bh14_uid164_Out0(1);
   bh14_w85_5 <= Compressor_6_3_F50_uid99_bh14_uid164_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid166_In0 <= "" & bh14_w84_0 & bh14_w84_1 & bh14_w84_2 & bh14_w84_3;
   Compressor_14_3_F50_uid63_bh14_uid166_In1 <= "" & bh14_w85_0;
   Compressor_14_3_F50_uid63_uid166: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid166_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid166_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid166_Out0_copy167);
   Compressor_14_3_F50_uid63_bh14_uid166_Out0 <= Compressor_14_3_F50_uid63_bh14_uid166_Out0_copy167; -- output copy to hold a pipeline register if needed

   bh14_w84_7 <= Compressor_14_3_F50_uid63_bh14_uid166_Out0(0);
   bh14_w85_6 <= Compressor_14_3_F50_uid63_bh14_uid166_Out0(1);
   bh14_w86_5 <= Compressor_14_3_F50_uid63_bh14_uid166_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid168_In0 <= "" & bh14_w85_1 & bh14_w85_2 & bh14_w85_3 & bh14_w85_4;
   Compressor_14_3_F50_uid63_bh14_uid168_In1 <= "" & bh14_w86_0;
   Compressor_14_3_F50_uid63_uid168: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid168_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid168_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid168_Out0_copy169);
   Compressor_14_3_F50_uid63_bh14_uid168_Out0 <= Compressor_14_3_F50_uid63_bh14_uid168_Out0_copy169; -- output copy to hold a pipeline register if needed

   bh14_w85_7 <= Compressor_14_3_F50_uid63_bh14_uid168_Out0(0);
   bh14_w86_6 <= Compressor_14_3_F50_uid63_bh14_uid168_Out0(1);
   bh14_w87_5 <= Compressor_14_3_F50_uid63_bh14_uid168_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid170_In0 <= "" & bh14_w86_1 & bh14_w86_2 & bh14_w86_3 & bh14_w86_4;
   Compressor_14_3_F50_uid63_bh14_uid170_In1 <= "" & bh14_w87_0;
   Compressor_14_3_F50_uid63_uid170: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid170_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid170_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid170_Out0_copy171);
   Compressor_14_3_F50_uid63_bh14_uid170_Out0 <= Compressor_14_3_F50_uid63_bh14_uid170_Out0_copy171; -- output copy to hold a pipeline register if needed

   bh14_w86_7 <= Compressor_14_3_F50_uid63_bh14_uid170_Out0(0);
   bh14_w87_6 <= Compressor_14_3_F50_uid63_bh14_uid170_Out0(1);
   bh14_w88_5 <= Compressor_14_3_F50_uid63_bh14_uid170_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid172_In0 <= "" & bh14_w87_1 & bh14_w87_2 & bh14_w87_3 & bh14_w87_4;
   Compressor_14_3_F50_uid63_bh14_uid172_In1 <= "" & bh14_w88_0;
   Compressor_14_3_F50_uid63_uid172: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid172_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid172_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid172_Out0_copy173);
   Compressor_14_3_F50_uid63_bh14_uid172_Out0 <= Compressor_14_3_F50_uid63_bh14_uid172_Out0_copy173; -- output copy to hold a pipeline register if needed

   bh14_w87_7 <= Compressor_14_3_F50_uid63_bh14_uid172_Out0(0);
   bh14_w88_6 <= Compressor_14_3_F50_uid63_bh14_uid172_Out0(1);
   bh14_w89_5 <= Compressor_14_3_F50_uid63_bh14_uid172_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid174_In0 <= "" & bh14_w88_1 & bh14_w88_2 & bh14_w88_3 & bh14_w88_4;
   Compressor_14_3_F50_uid63_bh14_uid174_In1 <= "" & bh14_w89_0;
   Compressor_14_3_F50_uid63_uid174: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid174_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid174_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid174_Out0_copy175);
   Compressor_14_3_F50_uid63_bh14_uid174_Out0 <= Compressor_14_3_F50_uid63_bh14_uid174_Out0_copy175; -- output copy to hold a pipeline register if needed

   bh14_w88_7 <= Compressor_14_3_F50_uid63_bh14_uid174_Out0(0);
   bh14_w89_6 <= Compressor_14_3_F50_uid63_bh14_uid174_Out0(1);
   bh14_w90_5 <= Compressor_14_3_F50_uid63_bh14_uid174_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid176_In0 <= "" & bh14_w89_1 & bh14_w89_2 & bh14_w89_3 & bh14_w89_4;
   Compressor_14_3_F50_uid63_bh14_uid176_In1 <= "" & bh14_w90_0;
   Compressor_14_3_F50_uid63_uid176: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid176_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid176_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid176_Out0_copy177);
   Compressor_14_3_F50_uid63_bh14_uid176_Out0 <= Compressor_14_3_F50_uid63_bh14_uid176_Out0_copy177; -- output copy to hold a pipeline register if needed

   bh14_w89_7 <= Compressor_14_3_F50_uid63_bh14_uid176_Out0(0);
   bh14_w90_6 <= Compressor_14_3_F50_uid63_bh14_uid176_Out0(1);
   bh14_w91_5 <= Compressor_14_3_F50_uid63_bh14_uid176_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid178_In0 <= "" & bh14_w90_1 & bh14_w90_2 & bh14_w90_3 & bh14_w90_4;
   Compressor_14_3_F50_uid63_bh14_uid178_In1 <= "" & bh14_w91_0;
   Compressor_14_3_F50_uid63_uid178: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid178_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid178_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid178_Out0_copy179);
   Compressor_14_3_F50_uid63_bh14_uid178_Out0 <= Compressor_14_3_F50_uid63_bh14_uid178_Out0_copy179; -- output copy to hold a pipeline register if needed

   bh14_w90_7 <= Compressor_14_3_F50_uid63_bh14_uid178_Out0(0);
   bh14_w91_6 <= Compressor_14_3_F50_uid63_bh14_uid178_Out0(1);
   bh14_w92_5 <= Compressor_14_3_F50_uid63_bh14_uid178_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid180_In0 <= "" & bh14_w91_1 & bh14_w91_2 & bh14_w91_3 & bh14_w91_4;
   Compressor_14_3_F50_uid63_bh14_uid180_In1 <= "" & bh14_w92_0;
   Compressor_14_3_F50_uid63_uid180: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid180_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid180_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid180_Out0_copy181);
   Compressor_14_3_F50_uid63_bh14_uid180_Out0 <= Compressor_14_3_F50_uid63_bh14_uid180_Out0_copy181; -- output copy to hold a pipeline register if needed

   bh14_w91_7 <= Compressor_14_3_F50_uid63_bh14_uid180_Out0(0);
   bh14_w92_6 <= Compressor_14_3_F50_uid63_bh14_uid180_Out0(1);
   bh14_w93_5 <= Compressor_14_3_F50_uid63_bh14_uid180_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid182_In0 <= "" & bh14_w92_1 & bh14_w92_2 & bh14_w92_3 & bh14_w92_4;
   Compressor_14_3_F50_uid63_bh14_uid182_In1 <= "" & bh14_w93_0;
   Compressor_14_3_F50_uid63_uid182: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid182_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid182_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid182_Out0_copy183);
   Compressor_14_3_F50_uid63_bh14_uid182_Out0 <= Compressor_14_3_F50_uid63_bh14_uid182_Out0_copy183; -- output copy to hold a pipeline register if needed

   bh14_w92_7 <= Compressor_14_3_F50_uid63_bh14_uid182_Out0(0);
   bh14_w93_6 <= Compressor_14_3_F50_uid63_bh14_uid182_Out0(1);
   bh14_w94_4 <= Compressor_14_3_F50_uid63_bh14_uid182_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid184_In0 <= "" & bh14_w93_1 & bh14_w93_2 & bh14_w93_3 & bh14_w93_4;
   Compressor_14_3_F50_uid63_bh14_uid184_In1 <= "" & bh14_w94_0;
   Compressor_14_3_F50_uid63_uid184: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid184_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid184_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid184_Out0_copy185);
   Compressor_14_3_F50_uid63_bh14_uid184_Out0 <= Compressor_14_3_F50_uid63_bh14_uid184_Out0_copy185; -- output copy to hold a pipeline register if needed

   bh14_w93_7 <= Compressor_14_3_F50_uid63_bh14_uid184_Out0(0);
   bh14_w94_5 <= Compressor_14_3_F50_uid63_bh14_uid184_Out0(1);
   bh14_w95_4 <= Compressor_14_3_F50_uid63_bh14_uid184_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid186_In0 <= "" & bh14_w94_1 & bh14_w94_2 & bh14_w94_3;
   Compressor_3_2_F50_uid49_uid186: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid186_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid186_Out0_copy187);
   Compressor_3_2_F50_uid49_bh14_uid186_Out0 <= Compressor_3_2_F50_uid49_bh14_uid186_Out0_copy187; -- output copy to hold a pipeline register if needed

   bh14_w94_6 <= Compressor_3_2_F50_uid49_bh14_uid186_Out0(0);
   bh14_w95_5 <= Compressor_3_2_F50_uid49_bh14_uid186_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid188_In0 <= "" & bh14_w95_0 & bh14_w95_1 & bh14_w95_2 & bh14_w95_3;
   Compressor_14_3_F50_uid63_bh14_uid188_In1 <= "" & bh14_w96_0;
   Compressor_14_3_F50_uid63_uid188: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid188_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid188_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid188_Out0_copy189);
   Compressor_14_3_F50_uid63_bh14_uid188_Out0 <= Compressor_14_3_F50_uid63_bh14_uid188_Out0_copy189; -- output copy to hold a pipeline register if needed

   bh14_w95_6 <= Compressor_14_3_F50_uid63_bh14_uid188_Out0(0);
   bh14_w96_4 <= Compressor_14_3_F50_uid63_bh14_uid188_Out0(1);
   bh14_w97_4 <= Compressor_14_3_F50_uid63_bh14_uid188_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid190_In0 <= "" & bh14_w96_1 & bh14_w96_2 & bh14_w96_3;
   Compressor_3_2_F50_uid49_uid190: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid190_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid190_Out0_copy191);
   Compressor_3_2_F50_uid49_bh14_uid190_Out0 <= Compressor_3_2_F50_uid49_bh14_uid190_Out0_copy191; -- output copy to hold a pipeline register if needed

   bh14_w96_5 <= Compressor_3_2_F50_uid49_bh14_uid190_Out0(0);
   bh14_w97_5 <= Compressor_3_2_F50_uid49_bh14_uid190_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid192_In0 <= "" & bh14_w97_0 & bh14_w97_1 & bh14_w97_2 & bh14_w97_3;
   Compressor_14_3_F50_uid63_bh14_uid192_In1 <= "" & bh14_w98_0;
   Compressor_14_3_F50_uid63_uid192: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid192_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid192_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid192_Out0_copy193);
   Compressor_14_3_F50_uid63_bh14_uid192_Out0 <= Compressor_14_3_F50_uid63_bh14_uid192_Out0_copy193; -- output copy to hold a pipeline register if needed

   bh14_w97_6 <= Compressor_14_3_F50_uid63_bh14_uid192_Out0(0);
   bh14_w98_4 <= Compressor_14_3_F50_uid63_bh14_uid192_Out0(1);
   bh14_w99_4 <= Compressor_14_3_F50_uid63_bh14_uid192_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid194_In0 <= "" & bh14_w98_1 & bh14_w98_2 & bh14_w98_3;
   Compressor_3_2_F50_uid49_uid194: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid194_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid194_Out0_copy195);
   Compressor_3_2_F50_uid49_bh14_uid194_Out0 <= Compressor_3_2_F50_uid49_bh14_uid194_Out0_copy195; -- output copy to hold a pipeline register if needed

   bh14_w98_5 <= Compressor_3_2_F50_uid49_bh14_uid194_Out0(0);
   bh14_w99_5 <= Compressor_3_2_F50_uid49_bh14_uid194_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid196_In0 <= "" & bh14_w99_0 & bh14_w99_1 & bh14_w99_2 & bh14_w99_3;
   Compressor_14_3_F50_uid63_bh14_uid196_In1 <= "" & bh14_w100_0;
   Compressor_14_3_F50_uid63_uid196: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid196_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid196_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid196_Out0_copy197);
   Compressor_14_3_F50_uid63_bh14_uid196_Out0 <= Compressor_14_3_F50_uid63_bh14_uid196_Out0_copy197; -- output copy to hold a pipeline register if needed

   bh14_w99_6 <= Compressor_14_3_F50_uid63_bh14_uid196_Out0(0);
   bh14_w100_4 <= Compressor_14_3_F50_uid63_bh14_uid196_Out0(1);
   bh14_w101_4 <= Compressor_14_3_F50_uid63_bh14_uid196_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid198_In0 <= "" & bh14_w100_1 & bh14_w100_2 & bh14_w100_3;
   Compressor_3_2_F50_uid49_uid198: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid198_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid198_Out0_copy199);
   Compressor_3_2_F50_uid49_bh14_uid198_Out0 <= Compressor_3_2_F50_uid49_bh14_uid198_Out0_copy199; -- output copy to hold a pipeline register if needed

   bh14_w100_5 <= Compressor_3_2_F50_uid49_bh14_uid198_Out0(0);
   bh14_w101_5 <= Compressor_3_2_F50_uid49_bh14_uid198_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid200_In0 <= "" & bh14_w101_0 & bh14_w101_1 & bh14_w101_2 & bh14_w101_3;
   Compressor_14_3_F50_uid63_bh14_uid200_In1 <= "" & bh14_w102_0;
   Compressor_14_3_F50_uid63_uid200: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid200_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid200_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid200_Out0_copy201);
   Compressor_14_3_F50_uid63_bh14_uid200_Out0 <= Compressor_14_3_F50_uid63_bh14_uid200_Out0_copy201; -- output copy to hold a pipeline register if needed

   bh14_w101_6 <= Compressor_14_3_F50_uid63_bh14_uid200_Out0(0);
   bh14_w102_4 <= Compressor_14_3_F50_uid63_bh14_uid200_Out0(1);
   bh14_w103_4 <= Compressor_14_3_F50_uid63_bh14_uid200_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid202_In0 <= "" & bh14_w102_1 & bh14_w102_2 & bh14_w102_3;
   Compressor_3_2_F50_uid49_uid202: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid202_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid202_Out0_copy203);
   Compressor_3_2_F50_uid49_bh14_uid202_Out0 <= Compressor_3_2_F50_uid49_bh14_uid202_Out0_copy203; -- output copy to hold a pipeline register if needed

   bh14_w102_5 <= Compressor_3_2_F50_uid49_bh14_uid202_Out0(0);
   bh14_w103_5 <= Compressor_3_2_F50_uid49_bh14_uid202_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid204_In0 <= "" & bh14_w103_0 & bh14_w103_1 & bh14_w103_2 & bh14_w103_3;
   Compressor_14_3_F50_uid63_bh14_uid204_In1 <= "" & bh14_w104_0;
   Compressor_14_3_F50_uid63_uid204: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid204_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid204_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid204_Out0_copy205);
   Compressor_14_3_F50_uid63_bh14_uid204_Out0 <= Compressor_14_3_F50_uid63_bh14_uid204_Out0_copy205; -- output copy to hold a pipeline register if needed

   bh14_w103_6 <= Compressor_14_3_F50_uid63_bh14_uid204_Out0(0);
   bh14_w104_4 <= Compressor_14_3_F50_uid63_bh14_uid204_Out0(1);
   bh14_w105_4 <= Compressor_14_3_F50_uid63_bh14_uid204_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid206_In0 <= "" & bh14_w104_1 & bh14_w104_2 & bh14_w104_3;
   Compressor_3_2_F50_uid49_uid206: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid206_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid206_Out0_copy207);
   Compressor_3_2_F50_uid49_bh14_uid206_Out0 <= Compressor_3_2_F50_uid49_bh14_uid206_Out0_copy207; -- output copy to hold a pipeline register if needed

   bh14_w104_5 <= Compressor_3_2_F50_uid49_bh14_uid206_Out0(0);
   bh14_w105_5 <= Compressor_3_2_F50_uid49_bh14_uid206_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid208_In0 <= "" & bh14_w105_0 & bh14_w105_1 & bh14_w105_2 & bh14_w105_3;
   Compressor_14_3_F50_uid63_bh14_uid208_In1 <= "" & bh14_w106_0;
   Compressor_14_3_F50_uid63_uid208: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid208_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid208_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid208_Out0_copy209);
   Compressor_14_3_F50_uid63_bh14_uid208_Out0 <= Compressor_14_3_F50_uid63_bh14_uid208_Out0_copy209; -- output copy to hold a pipeline register if needed

   bh14_w105_6 <= Compressor_14_3_F50_uid63_bh14_uid208_Out0(0);
   bh14_w106_4 <= Compressor_14_3_F50_uid63_bh14_uid208_Out0(1);
   bh14_w107_4 <= Compressor_14_3_F50_uid63_bh14_uid208_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid210_In0 <= "" & bh14_w106_1 & bh14_w106_2 & bh14_w106_3;
   Compressor_3_2_F50_uid49_uid210: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid210_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid210_Out0_copy211);
   Compressor_3_2_F50_uid49_bh14_uid210_Out0 <= Compressor_3_2_F50_uid49_bh14_uid210_Out0_copy211; -- output copy to hold a pipeline register if needed

   bh14_w106_5 <= Compressor_3_2_F50_uid49_bh14_uid210_Out0(0);
   bh14_w107_5 <= Compressor_3_2_F50_uid49_bh14_uid210_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid212_In0 <= "" & bh14_w107_0 & bh14_w107_1 & bh14_w107_2 & bh14_w107_3;
   Compressor_14_3_F50_uid63_bh14_uid212_In1 <= "" & "0";
   Compressor_14_3_F50_uid63_uid212: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid212_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid212_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid212_Out0_copy213);
   Compressor_14_3_F50_uid63_bh14_uid212_Out0 <= Compressor_14_3_F50_uid63_bh14_uid212_Out0_copy213; -- output copy to hold a pipeline register if needed

   bh14_w107_6 <= Compressor_14_3_F50_uid63_bh14_uid212_Out0(0);
   bh14_w108_3 <= Compressor_14_3_F50_uid63_bh14_uid212_Out0(1);
   bh14_w109_3 <= Compressor_14_3_F50_uid63_bh14_uid212_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid214_In0 <= "" & bh14_w108_0 & bh14_w108_1 & bh14_w108_2;
   Compressor_3_2_F50_uid49_uid214: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid214_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid214_Out0_copy215);
   Compressor_3_2_F50_uid49_bh14_uid214_Out0 <= Compressor_3_2_F50_uid49_bh14_uid214_Out0_copy215; -- output copy to hold a pipeline register if needed

   bh14_w108_4 <= Compressor_3_2_F50_uid49_bh14_uid214_Out0(0);
   bh14_w109_4 <= Compressor_3_2_F50_uid49_bh14_uid214_Out0(1);

   Compressor_23_3_F50_uid41_bh14_uid216_In0 <= "" & bh14_w109_0 & bh14_w109_1 & bh14_w109_2;
   Compressor_23_3_F50_uid41_bh14_uid216_In1 <= "" & bh14_w110_0 & bh14_w110_1;
   Compressor_23_3_F50_uid41_uid216: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid216_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid216_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid216_Out0_copy217);
   Compressor_23_3_F50_uid41_bh14_uid216_Out0 <= Compressor_23_3_F50_uid41_bh14_uid216_Out0_copy217; -- output copy to hold a pipeline register if needed

   bh14_w109_5 <= Compressor_23_3_F50_uid41_bh14_uid216_Out0(0);
   bh14_w110_3 <= Compressor_23_3_F50_uid41_bh14_uid216_Out0(1);
   bh14_w111_2 <= Compressor_23_3_F50_uid41_bh14_uid216_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid218_In0 <= "" & bh14_w111_0 & bh14_w111_1 & "0";
   Compressor_23_3_F50_uid41_bh14_uid218_In1 <= "" & bh14_w112_0 & bh14_w112_1;
   Compressor_23_3_F50_uid41_uid218: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid218_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid218_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid218_Out0_copy219);
   Compressor_23_3_F50_uid41_bh14_uid218_Out0 <= Compressor_23_3_F50_uid41_bh14_uid218_Out0_copy219; -- output copy to hold a pipeline register if needed

   bh14_w111_3 <= Compressor_23_3_F50_uid41_bh14_uid218_Out0(0);
   bh14_w112_2 <= Compressor_23_3_F50_uid41_bh14_uid218_Out0(1);
   bh14_w113_2 <= Compressor_23_3_F50_uid41_bh14_uid218_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid220_In0 <= "" & bh14_w113_0 & bh14_w113_1 & "0";
   Compressor_23_3_F50_uid41_bh14_uid220_In1 <= "" & bh14_w114_0 & bh14_w114_1;
   Compressor_23_3_F50_uid41_uid220: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid220_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid220_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid220_Out0_copy221);
   Compressor_23_3_F50_uid41_bh14_uid220_Out0 <= Compressor_23_3_F50_uid41_bh14_uid220_Out0_copy221; -- output copy to hold a pipeline register if needed

   bh14_w113_3 <= Compressor_23_3_F50_uid41_bh14_uid220_Out0(0);
   bh14_w114_2 <= Compressor_23_3_F50_uid41_bh14_uid220_Out0(1);
   bh14_w115_2 <= Compressor_23_3_F50_uid41_bh14_uid220_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid222_In0 <= "" & bh14_w115_0 & bh14_w115_1 & "0";
   Compressor_23_3_F50_uid41_bh14_uid222_In1 <= "" & bh14_w116_0 & bh14_w116_1;
   Compressor_23_3_F50_uid41_uid222: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid222_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid222_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid222_Out0_copy223);
   Compressor_23_3_F50_uid41_bh14_uid222_Out0 <= Compressor_23_3_F50_uid41_bh14_uid222_Out0_copy223; -- output copy to hold a pipeline register if needed

   bh14_w115_3 <= Compressor_23_3_F50_uid41_bh14_uid222_Out0(0);
   bh14_w116_2 <= Compressor_23_3_F50_uid41_bh14_uid222_Out0(1);
   bh14_w117_2 <= Compressor_23_3_F50_uid41_bh14_uid222_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid224_In0 <= "" & bh14_w117_0 & bh14_w117_1 & "0";
   Compressor_23_3_F50_uid41_bh14_uid224_In1 <= "" & bh14_w118_0 & bh14_w118_1;
   Compressor_23_3_F50_uid41_uid224: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid224_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid224_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid224_Out0_copy225);
   Compressor_23_3_F50_uid41_bh14_uid224_Out0 <= Compressor_23_3_F50_uid41_bh14_uid224_Out0_copy225; -- output copy to hold a pipeline register if needed

   bh14_w117_3 <= Compressor_23_3_F50_uid41_bh14_uid224_Out0(0);
   bh14_w118_2 <= Compressor_23_3_F50_uid41_bh14_uid224_Out0(1);
   bh14_w119_2 <= Compressor_23_3_F50_uid41_bh14_uid224_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid226_In0 <= "" & bh14_w119_0 & bh14_w119_1 & "0";
   Compressor_23_3_F50_uid41_bh14_uid226_In1 <= "" & bh14_w120_0 & bh14_w120_1;
   Compressor_23_3_F50_uid41_uid226: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid226_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid226_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid226_Out0_copy227);
   Compressor_23_3_F50_uid41_bh14_uid226_Out0 <= Compressor_23_3_F50_uid41_bh14_uid226_Out0_copy227; -- output copy to hold a pipeline register if needed

   bh14_w119_3 <= Compressor_23_3_F50_uid41_bh14_uid226_Out0(0);
   bh14_w120_2 <= Compressor_23_3_F50_uid41_bh14_uid226_Out0(1);
   bh14_w121_1 <= Compressor_23_3_F50_uid41_bh14_uid226_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid228_In0 <= "" & bh14_w19_3 & bh14_w19_2 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid228_In1 <= "" & bh14_w20_2;
   Compressor_14_3_F50_uid63_uid228: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid228_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid228_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid228_Out0_copy229);
   Compressor_14_3_F50_uid63_bh14_uid228_Out0 <= Compressor_14_3_F50_uid63_bh14_uid228_Out0_copy229; -- output copy to hold a pipeline register if needed

   bh14_w19_4 <= Compressor_14_3_F50_uid63_bh14_uid228_Out0(0);
   bh14_w20_3 <= Compressor_14_3_F50_uid63_bh14_uid228_Out0(1);
   bh14_w21_4 <= Compressor_14_3_F50_uid63_bh14_uid228_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid230_In0 <= "" & bh14_w21_3 & bh14_w21_2 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid230_In1 <= "" & bh14_w22_2;
   Compressor_14_3_F50_uid63_uid230: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid230_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid230_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid230_Out0_copy231);
   Compressor_14_3_F50_uid63_bh14_uid230_Out0 <= Compressor_14_3_F50_uid63_bh14_uid230_Out0_copy231; -- output copy to hold a pipeline register if needed

   bh14_w21_5 <= Compressor_14_3_F50_uid63_bh14_uid230_Out0(0);
   bh14_w22_3 <= Compressor_14_3_F50_uid63_bh14_uid230_Out0(1);
   bh14_w23_4 <= Compressor_14_3_F50_uid63_bh14_uid230_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid232_In0 <= "" & bh14_w23_3 & bh14_w23_2 & "0";
   Compressor_23_3_F50_uid41_bh14_uid232_In1 <= "" & bh14_w24_4 & bh14_w24_3;
   Compressor_23_3_F50_uid41_uid232: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid232_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid232_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid232_Out0_copy233);
   Compressor_23_3_F50_uid41_bh14_uid232_Out0 <= Compressor_23_3_F50_uid41_bh14_uid232_Out0_copy233; -- output copy to hold a pipeline register if needed

   bh14_w23_5 <= Compressor_23_3_F50_uid41_bh14_uid232_Out0(0);
   bh14_w24_5 <= Compressor_23_3_F50_uid41_bh14_uid232_Out0(1);
   bh14_w25_4 <= Compressor_23_3_F50_uid41_bh14_uid232_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid234_In0 <= "" & bh14_w25_3 & bh14_w25_2 & "0";
   Compressor_23_3_F50_uid41_bh14_uid234_In1 <= "" & bh14_w26_4 & bh14_w26_3;
   Compressor_23_3_F50_uid41_uid234: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid234_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid234_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid234_Out0_copy235);
   Compressor_23_3_F50_uid41_bh14_uid234_Out0 <= Compressor_23_3_F50_uid41_bh14_uid234_Out0_copy235; -- output copy to hold a pipeline register if needed

   bh14_w25_5 <= Compressor_23_3_F50_uid41_bh14_uid234_Out0(0);
   bh14_w26_5 <= Compressor_23_3_F50_uid41_bh14_uid234_Out0(1);
   bh14_w27_4 <= Compressor_23_3_F50_uid41_bh14_uid234_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid236_In0 <= "" & bh14_w27_3 & bh14_w27_2 & "0";
   Compressor_23_3_F50_uid41_bh14_uid236_In1 <= "" & bh14_w28_4 & bh14_w28_3;
   Compressor_23_3_F50_uid41_uid236: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid236_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid236_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid236_Out0_copy237);
   Compressor_23_3_F50_uid41_bh14_uid236_Out0 <= Compressor_23_3_F50_uid41_bh14_uid236_Out0_copy237; -- output copy to hold a pipeline register if needed

   bh14_w27_5 <= Compressor_23_3_F50_uid41_bh14_uid236_Out0(0);
   bh14_w28_5 <= Compressor_23_3_F50_uid41_bh14_uid236_Out0(1);
   bh14_w29_4 <= Compressor_23_3_F50_uid41_bh14_uid236_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid238_In0 <= "" & bh14_w29_3 & bh14_w29_2 & "0";
   Compressor_23_3_F50_uid41_bh14_uid238_In1 <= "" & bh14_w30_4 & bh14_w30_3;
   Compressor_23_3_F50_uid41_uid238: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid238_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid238_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid238_Out0_copy239);
   Compressor_23_3_F50_uid41_bh14_uid238_Out0 <= Compressor_23_3_F50_uid41_bh14_uid238_Out0_copy239; -- output copy to hold a pipeline register if needed

   bh14_w29_5 <= Compressor_23_3_F50_uid41_bh14_uid238_Out0(0);
   bh14_w30_5 <= Compressor_23_3_F50_uid41_bh14_uid238_Out0(1);
   bh14_w31_4 <= Compressor_23_3_F50_uid41_bh14_uid238_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid240_In0 <= "" & bh14_w31_3 & bh14_w31_2 & "0";
   Compressor_23_3_F50_uid41_bh14_uid240_In1 <= "" & bh14_w32_4 & bh14_w32_3;
   Compressor_23_3_F50_uid41_uid240: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid240_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid240_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid240_Out0_copy241);
   Compressor_23_3_F50_uid41_bh14_uid240_Out0 <= Compressor_23_3_F50_uid41_bh14_uid240_Out0_copy241; -- output copy to hold a pipeline register if needed

   bh14_w31_5 <= Compressor_23_3_F50_uid41_bh14_uid240_Out0(0);
   bh14_w32_5 <= Compressor_23_3_F50_uid41_bh14_uid240_Out0(1);
   bh14_w33_4 <= Compressor_23_3_F50_uid41_bh14_uid240_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid242_In0 <= "" & bh14_w33_3 & bh14_w33_2 & "0";
   Compressor_23_3_F50_uid41_bh14_uid242_In1 <= "" & bh14_w34_5 & bh14_w34_4;
   Compressor_23_3_F50_uid41_uid242: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid242_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid242_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid242_Out0_copy243);
   Compressor_23_3_F50_uid41_bh14_uid242_Out0 <= Compressor_23_3_F50_uid41_bh14_uid242_Out0_copy243; -- output copy to hold a pipeline register if needed

   bh14_w33_5 <= Compressor_23_3_F50_uid41_bh14_uid242_Out0(0);
   bh14_w34_6 <= Compressor_23_3_F50_uid41_bh14_uid242_Out0(1);
   bh14_w35_6 <= Compressor_23_3_F50_uid41_bh14_uid242_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid244_In0 <= "" & bh14_w35_5 & bh14_w35_4 & "0";
   Compressor_3_2_F50_uid49_uid244: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid244_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid244_Out0_copy245);
   Compressor_3_2_F50_uid49_bh14_uid244_Out0 <= Compressor_3_2_F50_uid49_bh14_uid244_Out0_copy245; -- output copy to hold a pipeline register if needed

   bh14_w35_7 <= Compressor_3_2_F50_uid49_bh14_uid244_Out0(0);
   bh14_w36_7 <= Compressor_3_2_F50_uid49_bh14_uid244_Out0(1);

   Compressor_23_3_F50_uid41_bh14_uid246_In0 <= "" & bh14_w36_6 & bh14_w36_5 & bh14_w36_4;
   Compressor_23_3_F50_uid41_bh14_uid246_In1 <= "" & bh14_w37_5 & bh14_w37_4;
   Compressor_23_3_F50_uid41_uid246: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid246_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid246_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid246_Out0_copy247);
   Compressor_23_3_F50_uid41_bh14_uid246_Out0 <= Compressor_23_3_F50_uid41_bh14_uid246_Out0_copy247; -- output copy to hold a pipeline register if needed

   bh14_w36_8 <= Compressor_23_3_F50_uid41_bh14_uid246_Out0(0);
   bh14_w37_6 <= Compressor_23_3_F50_uid41_bh14_uid246_Out0(1);
   bh14_w38_7 <= Compressor_23_3_F50_uid41_bh14_uid246_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid248_In0 <= "" & bh14_w38_6 & bh14_w38_5 & bh14_w38_4;
   Compressor_23_3_F50_uid41_bh14_uid248_In1 <= "" & bh14_w39_5 & bh14_w39_4;
   Compressor_23_3_F50_uid41_uid248: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid248_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid248_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid248_Out0_copy249);
   Compressor_23_3_F50_uid41_bh14_uid248_Out0 <= Compressor_23_3_F50_uid41_bh14_uid248_Out0_copy249; -- output copy to hold a pipeline register if needed

   bh14_w38_8 <= Compressor_23_3_F50_uid41_bh14_uid248_Out0(0);
   bh14_w39_6 <= Compressor_23_3_F50_uid41_bh14_uid248_Out0(1);
   bh14_w40_7 <= Compressor_23_3_F50_uid41_bh14_uid248_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid250_In0 <= "" & bh14_w40_6 & bh14_w40_5 & bh14_w40_4;
   Compressor_23_3_F50_uid41_bh14_uid250_In1 <= "" & bh14_w41_5 & bh14_w41_4;
   Compressor_23_3_F50_uid41_uid250: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid250_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid250_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid250_Out0_copy251);
   Compressor_23_3_F50_uid41_bh14_uid250_Out0 <= Compressor_23_3_F50_uid41_bh14_uid250_Out0_copy251; -- output copy to hold a pipeline register if needed

   bh14_w40_8 <= Compressor_23_3_F50_uid41_bh14_uid250_Out0(0);
   bh14_w41_6 <= Compressor_23_3_F50_uid41_bh14_uid250_Out0(1);
   bh14_w42_7 <= Compressor_23_3_F50_uid41_bh14_uid250_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid252_In0 <= "" & bh14_w42_6 & bh14_w42_5 & bh14_w42_4;
   Compressor_23_3_F50_uid41_bh14_uid252_In1 <= "" & bh14_w43_5 & bh14_w43_4;
   Compressor_23_3_F50_uid41_uid252: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid252_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid252_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid252_Out0_copy253);
   Compressor_23_3_F50_uid41_bh14_uid252_Out0 <= Compressor_23_3_F50_uid41_bh14_uid252_Out0_copy253; -- output copy to hold a pipeline register if needed

   bh14_w42_8 <= Compressor_23_3_F50_uid41_bh14_uid252_Out0(0);
   bh14_w43_6 <= Compressor_23_3_F50_uid41_bh14_uid252_Out0(1);
   bh14_w44_7 <= Compressor_23_3_F50_uid41_bh14_uid252_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid254_In0 <= "" & bh14_w44_6 & bh14_w44_5 & bh14_w44_4;
   Compressor_23_3_F50_uid41_bh14_uid254_In1 <= "" & bh14_w45_5 & bh14_w45_4;
   Compressor_23_3_F50_uid41_uid254: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid254_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid254_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid254_Out0_copy255);
   Compressor_23_3_F50_uid41_bh14_uid254_Out0 <= Compressor_23_3_F50_uid41_bh14_uid254_Out0_copy255; -- output copy to hold a pipeline register if needed

   bh14_w44_8 <= Compressor_23_3_F50_uid41_bh14_uid254_Out0(0);
   bh14_w45_6 <= Compressor_23_3_F50_uid41_bh14_uid254_Out0(1);
   bh14_w46_7 <= Compressor_23_3_F50_uid41_bh14_uid254_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid256_In0 <= "" & bh14_w46_6 & bh14_w46_5 & bh14_w46_4;
   Compressor_23_3_F50_uid41_bh14_uid256_In1 <= "" & bh14_w47_5 & bh14_w47_4;
   Compressor_23_3_F50_uid41_uid256: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid256_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid256_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid256_Out0_copy257);
   Compressor_23_3_F50_uid41_bh14_uid256_Out0 <= Compressor_23_3_F50_uid41_bh14_uid256_Out0_copy257; -- output copy to hold a pipeline register if needed

   bh14_w46_8 <= Compressor_23_3_F50_uid41_bh14_uid256_Out0(0);
   bh14_w47_6 <= Compressor_23_3_F50_uid41_bh14_uid256_Out0(1);
   bh14_w48_8 <= Compressor_23_3_F50_uid41_bh14_uid256_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid258_In0 <= "" & bh14_w48_7 & bh14_w48_6 & bh14_w48_5 & bh14_w48_4;
   Compressor_14_3_F50_uid63_bh14_uid258_In1 <= "" & bh14_w49_6;
   Compressor_14_3_F50_uid63_uid258: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid258_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid258_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid258_Out0_copy259);
   Compressor_14_3_F50_uid63_bh14_uid258_Out0 <= Compressor_14_3_F50_uid63_bh14_uid258_Out0_copy259; -- output copy to hold a pipeline register if needed

   bh14_w48_9 <= Compressor_14_3_F50_uid63_bh14_uid258_Out0(0);
   bh14_w49_7 <= Compressor_14_3_F50_uid63_bh14_uid258_Out0(1);
   bh14_w50_8 <= Compressor_14_3_F50_uid63_bh14_uid258_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid260_In0 <= "" & bh14_w50_7 & bh14_w50_6 & bh14_w50_5 & bh14_w50_4;
   Compressor_14_3_F50_uid63_bh14_uid260_In1 <= "" & "0";
   Compressor_14_3_F50_uid63_uid260: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid260_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid260_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid260_Out0_copy261);
   Compressor_14_3_F50_uid63_bh14_uid260_Out0 <= Compressor_14_3_F50_uid63_bh14_uid260_Out0_copy261; -- output copy to hold a pipeline register if needed

   bh14_w50_9 <= Compressor_14_3_F50_uid63_bh14_uid260_Out0(0);
   bh14_w51_9 <= Compressor_14_3_F50_uid63_bh14_uid260_Out0(1);
   bh14_w52_8 <= Compressor_14_3_F50_uid63_bh14_uid260_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid262_In0 <= "" & bh14_w51_8 & bh14_w51_7 & bh14_w51_6;
   Compressor_23_3_F50_uid41_bh14_uid262_In1 <= "" & bh14_w52_7 & bh14_w52_6;
   Compressor_23_3_F50_uid41_uid262: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid262_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid262_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid262_Out0_copy263);
   Compressor_23_3_F50_uid41_bh14_uid262_Out0 <= Compressor_23_3_F50_uid41_bh14_uid262_Out0_copy263; -- output copy to hold a pipeline register if needed

   bh14_w51_10 <= Compressor_23_3_F50_uid41_bh14_uid262_Out0(0);
   bh14_w52_9 <= Compressor_23_3_F50_uid41_bh14_uid262_Out0(1);
   bh14_w53_9 <= Compressor_23_3_F50_uid41_bh14_uid262_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid264_In0 <= "" & bh14_w53_8 & bh14_w53_7 & bh14_w53_6;
   Compressor_23_3_F50_uid41_bh14_uid264_In1 <= "" & bh14_w54_8 & bh14_w54_7;
   Compressor_23_3_F50_uid41_uid264: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid264_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid264_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid264_Out0_copy265);
   Compressor_23_3_F50_uid41_bh14_uid264_Out0 <= Compressor_23_3_F50_uid41_bh14_uid264_Out0_copy265; -- output copy to hold a pipeline register if needed

   bh14_w53_10 <= Compressor_23_3_F50_uid41_bh14_uid264_Out0(0);
   bh14_w54_9 <= Compressor_23_3_F50_uid41_bh14_uid264_Out0(1);
   bh14_w55_9 <= Compressor_23_3_F50_uid41_bh14_uid264_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid266_In0 <= "" & bh14_w55_8 & bh14_w55_7 & bh14_w55_6;
   Compressor_23_3_F50_uid41_bh14_uid266_In1 <= "" & bh14_w56_8 & bh14_w56_7;
   Compressor_23_3_F50_uid41_uid266: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid266_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid266_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid266_Out0_copy267);
   Compressor_23_3_F50_uid41_bh14_uid266_Out0 <= Compressor_23_3_F50_uid41_bh14_uid266_Out0_copy267; -- output copy to hold a pipeline register if needed

   bh14_w55_10 <= Compressor_23_3_F50_uid41_bh14_uid266_Out0(0);
   bh14_w56_9 <= Compressor_23_3_F50_uid41_bh14_uid266_Out0(1);
   bh14_w57_9 <= Compressor_23_3_F50_uid41_bh14_uid266_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid268_In0 <= "" & bh14_w57_8 & bh14_w57_7 & bh14_w57_6;
   Compressor_23_3_F50_uid41_bh14_uid268_In1 <= "" & bh14_w58_8 & bh14_w58_7;
   Compressor_23_3_F50_uid41_uid268: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid268_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid268_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid268_Out0_copy269);
   Compressor_23_3_F50_uid41_bh14_uid268_Out0 <= Compressor_23_3_F50_uid41_bh14_uid268_Out0_copy269; -- output copy to hold a pipeline register if needed

   bh14_w57_10 <= Compressor_23_3_F50_uid41_bh14_uid268_Out0(0);
   bh14_w58_9 <= Compressor_23_3_F50_uid41_bh14_uid268_Out0(1);
   bh14_w59_9 <= Compressor_23_3_F50_uid41_bh14_uid268_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid270_In0 <= "" & bh14_w59_8 & bh14_w59_7 & bh14_w59_6;
   Compressor_23_3_F50_uid41_bh14_uid270_In1 <= "" & bh14_w60_8 & bh14_w60_7;
   Compressor_23_3_F50_uid41_uid270: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid270_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid270_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid270_Out0_copy271);
   Compressor_23_3_F50_uid41_bh14_uid270_Out0 <= Compressor_23_3_F50_uid41_bh14_uid270_Out0_copy271; -- output copy to hold a pipeline register if needed

   bh14_w59_10 <= Compressor_23_3_F50_uid41_bh14_uid270_Out0(0);
   bh14_w60_9 <= Compressor_23_3_F50_uid41_bh14_uid270_Out0(1);
   bh14_w61_9 <= Compressor_23_3_F50_uid41_bh14_uid270_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid272_In0 <= "" & bh14_w61_8 & bh14_w61_7 & bh14_w61_6;
   Compressor_23_3_F50_uid41_bh14_uid272_In1 <= "" & bh14_w62_8 & bh14_w62_7;
   Compressor_23_3_F50_uid41_uid272: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid272_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid272_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid272_Out0_copy273);
   Compressor_23_3_F50_uid41_bh14_uid272_Out0 <= Compressor_23_3_F50_uid41_bh14_uid272_Out0_copy273; -- output copy to hold a pipeline register if needed

   bh14_w61_10 <= Compressor_23_3_F50_uid41_bh14_uid272_Out0(0);
   bh14_w62_9 <= Compressor_23_3_F50_uid41_bh14_uid272_Out0(1);
   bh14_w63_9 <= Compressor_23_3_F50_uid41_bh14_uid272_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid274_In0 <= "" & bh14_w63_8 & bh14_w63_7 & bh14_w63_6;
   Compressor_23_3_F50_uid41_bh14_uid274_In1 <= "" & bh14_w64_8 & bh14_w64_7;
   Compressor_23_3_F50_uid41_uid274: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid274_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid274_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid274_Out0_copy275);
   Compressor_23_3_F50_uid41_bh14_uid274_Out0 <= Compressor_23_3_F50_uid41_bh14_uid274_Out0_copy275; -- output copy to hold a pipeline register if needed

   bh14_w63_10 <= Compressor_23_3_F50_uid41_bh14_uid274_Out0(0);
   bh14_w64_9 <= Compressor_23_3_F50_uid41_bh14_uid274_Out0(1);
   bh14_w65_9 <= Compressor_23_3_F50_uid41_bh14_uid274_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid276_In0 <= "" & bh14_w65_8 & bh14_w65_7 & bh14_w65_6;
   Compressor_23_3_F50_uid41_bh14_uid276_In1 <= "" & bh14_w66_8 & bh14_w66_7;
   Compressor_23_3_F50_uid41_uid276: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid276_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid276_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid276_Out0_copy277);
   Compressor_23_3_F50_uid41_bh14_uid276_Out0 <= Compressor_23_3_F50_uid41_bh14_uid276_Out0_copy277; -- output copy to hold a pipeline register if needed

   bh14_w65_10 <= Compressor_23_3_F50_uid41_bh14_uid276_Out0(0);
   bh14_w66_9 <= Compressor_23_3_F50_uid41_bh14_uid276_Out0(1);
   bh14_w67_9 <= Compressor_23_3_F50_uid41_bh14_uid276_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid278_In0 <= "" & bh14_w67_8 & bh14_w67_7 & bh14_w67_6;
   Compressor_23_3_F50_uid41_bh14_uid278_In1 <= "" & bh14_w68_8 & bh14_w68_7;
   Compressor_23_3_F50_uid41_uid278: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid278_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid278_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid278_Out0_copy279);
   Compressor_23_3_F50_uid41_bh14_uid278_Out0 <= Compressor_23_3_F50_uid41_bh14_uid278_Out0_copy279; -- output copy to hold a pipeline register if needed

   bh14_w67_10 <= Compressor_23_3_F50_uid41_bh14_uid278_Out0(0);
   bh14_w68_9 <= Compressor_23_3_F50_uid41_bh14_uid278_Out0(1);
   bh14_w69_9 <= Compressor_23_3_F50_uid41_bh14_uid278_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid280_In0 <= "" & bh14_w69_8 & bh14_w69_7 & bh14_w69_6;
   Compressor_23_3_F50_uid41_bh14_uid280_In1 <= "" & bh14_w70_8 & bh14_w70_7;
   Compressor_23_3_F50_uid41_uid280: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid280_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid280_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid280_Out0_copy281);
   Compressor_23_3_F50_uid41_bh14_uid280_Out0 <= Compressor_23_3_F50_uid41_bh14_uid280_Out0_copy281; -- output copy to hold a pipeline register if needed

   bh14_w69_10 <= Compressor_23_3_F50_uid41_bh14_uid280_Out0(0);
   bh14_w70_9 <= Compressor_23_3_F50_uid41_bh14_uid280_Out0(1);
   bh14_w71_9 <= Compressor_23_3_F50_uid41_bh14_uid280_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid282_In0 <= "" & bh14_w71_8 & bh14_w71_7 & bh14_w71_6;
   Compressor_23_3_F50_uid41_bh14_uid282_In1 <= "" & bh14_w72_8 & bh14_w72_7;
   Compressor_23_3_F50_uid41_uid282: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid282_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid282_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid282_Out0_copy283);
   Compressor_23_3_F50_uid41_bh14_uid282_Out0 <= Compressor_23_3_F50_uid41_bh14_uid282_Out0_copy283; -- output copy to hold a pipeline register if needed

   bh14_w71_10 <= Compressor_23_3_F50_uid41_bh14_uid282_Out0(0);
   bh14_w72_9 <= Compressor_23_3_F50_uid41_bh14_uid282_Out0(1);
   bh14_w73_9 <= Compressor_23_3_F50_uid41_bh14_uid282_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid284_In0 <= "" & bh14_w73_8 & bh14_w73_7 & bh14_w73_6;
   Compressor_23_3_F50_uid41_bh14_uid284_In1 <= "" & bh14_w74_8 & bh14_w74_7;
   Compressor_23_3_F50_uid41_uid284: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid284_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid284_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid284_Out0_copy285);
   Compressor_23_3_F50_uid41_bh14_uid284_Out0 <= Compressor_23_3_F50_uid41_bh14_uid284_Out0_copy285; -- output copy to hold a pipeline register if needed

   bh14_w73_10 <= Compressor_23_3_F50_uid41_bh14_uid284_Out0(0);
   bh14_w74_9 <= Compressor_23_3_F50_uid41_bh14_uid284_Out0(1);
   bh14_w75_9 <= Compressor_23_3_F50_uid41_bh14_uid284_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid286_In0 <= "" & bh14_w75_8 & bh14_w75_7 & bh14_w75_6;
   Compressor_23_3_F50_uid41_bh14_uid286_In1 <= "" & bh14_w76_8 & bh14_w76_7;
   Compressor_23_3_F50_uid41_uid286: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid286_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid286_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid286_Out0_copy287);
   Compressor_23_3_F50_uid41_bh14_uid286_Out0 <= Compressor_23_3_F50_uid41_bh14_uid286_Out0_copy287; -- output copy to hold a pipeline register if needed

   bh14_w75_10 <= Compressor_23_3_F50_uid41_bh14_uid286_Out0(0);
   bh14_w76_9 <= Compressor_23_3_F50_uid41_bh14_uid286_Out0(1);
   bh14_w77_10 <= Compressor_23_3_F50_uid41_bh14_uid286_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid288_In0 <= "" & bh14_w77_9 & bh14_w77_8 & bh14_w77_7 & bh14_w77_6;
   Compressor_14_3_F50_uid63_bh14_uid288_In1 <= "" & "0";
   Compressor_14_3_F50_uid63_uid288: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid288_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid288_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid288_Out0_copy289);
   Compressor_14_3_F50_uid63_bh14_uid288_Out0 <= Compressor_14_3_F50_uid63_bh14_uid288_Out0_copy289; -- output copy to hold a pipeline register if needed

   bh14_w77_11 <= Compressor_14_3_F50_uid63_bh14_uid288_Out0(0);
   bh14_w78_9 <= Compressor_14_3_F50_uid63_bh14_uid288_Out0(1);
   bh14_w79_9 <= Compressor_14_3_F50_uid63_bh14_uid288_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid290_In0 <= "" & bh14_w78_8 & bh14_w78_7 & bh14_w78_6;
   Compressor_3_2_F50_uid49_uid290: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid290_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid290_Out0_copy291);
   Compressor_3_2_F50_uid49_bh14_uid290_Out0 <= Compressor_3_2_F50_uid49_bh14_uid290_Out0_copy291; -- output copy to hold a pipeline register if needed

   bh14_w78_10 <= Compressor_3_2_F50_uid49_bh14_uid290_Out0(0);
   bh14_w79_10 <= Compressor_3_2_F50_uid49_bh14_uid290_Out0(1);

   Compressor_23_3_F50_uid41_bh14_uid292_In0 <= "" & bh14_w79_8 & bh14_w79_7 & bh14_w79_6;
   Compressor_23_3_F50_uid41_bh14_uid292_In1 <= "" & bh14_w80_8 & bh14_w80_7;
   Compressor_23_3_F50_uid41_uid292: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid292_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid292_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid292_Out0_copy293);
   Compressor_23_3_F50_uid41_bh14_uid292_Out0 <= Compressor_23_3_F50_uid41_bh14_uid292_Out0_copy293; -- output copy to hold a pipeline register if needed

   bh14_w79_11 <= Compressor_23_3_F50_uid41_bh14_uid292_Out0(0);
   bh14_w80_9 <= Compressor_23_3_F50_uid41_bh14_uid292_Out0(1);
   bh14_w81_9 <= Compressor_23_3_F50_uid41_bh14_uid292_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid294_In0 <= "" & bh14_w81_8 & bh14_w81_7 & bh14_w81_6;
   Compressor_23_3_F50_uid41_bh14_uid294_In1 <= "" & bh14_w82_8 & bh14_w82_7;
   Compressor_23_3_F50_uid41_uid294: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid294_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid294_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid294_Out0_copy295);
   Compressor_23_3_F50_uid41_bh14_uid294_Out0 <= Compressor_23_3_F50_uid41_bh14_uid294_Out0_copy295; -- output copy to hold a pipeline register if needed

   bh14_w81_10 <= Compressor_23_3_F50_uid41_bh14_uid294_Out0(0);
   bh14_w82_9 <= Compressor_23_3_F50_uid41_bh14_uid294_Out0(1);
   bh14_w83_9 <= Compressor_23_3_F50_uid41_bh14_uid294_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid296_In0 <= "" & bh14_w83_8 & bh14_w83_7 & bh14_w83_6;
   Compressor_3_2_F50_uid49_uid296: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid296_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid296_Out0_copy297);
   Compressor_3_2_F50_uid49_bh14_uid296_Out0 <= Compressor_3_2_F50_uid49_bh14_uid296_Out0_copy297; -- output copy to hold a pipeline register if needed

   bh14_w83_10 <= Compressor_3_2_F50_uid49_bh14_uid296_Out0(0);
   bh14_w84_8 <= Compressor_3_2_F50_uid49_bh14_uid296_Out0(1);

   Compressor_14_3_F50_uid63_bh14_uid298_In0 <= "" & bh14_w84_7 & bh14_w84_6 & bh14_w84_5 & bh14_w84_4;
   Compressor_14_3_F50_uid63_bh14_uid298_In1 <= "" & "0";
   Compressor_14_3_F50_uid63_uid298: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid298_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid298_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid298_Out0_copy299);
   Compressor_14_3_F50_uid63_bh14_uid298_Out0 <= Compressor_14_3_F50_uid63_bh14_uid298_Out0_copy299; -- output copy to hold a pipeline register if needed

   bh14_w84_9 <= Compressor_14_3_F50_uid63_bh14_uid298_Out0(0);
   bh14_w85_8 <= Compressor_14_3_F50_uid63_bh14_uid298_Out0(1);
   bh14_w86_8 <= Compressor_14_3_F50_uid63_bh14_uid298_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid300_In0 <= "" & bh14_w85_7 & bh14_w85_6 & bh14_w85_5;
   Compressor_3_2_F50_uid49_uid300: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid300_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid300_Out0_copy301);
   Compressor_3_2_F50_uid49_bh14_uid300_Out0 <= Compressor_3_2_F50_uid49_bh14_uid300_Out0_copy301; -- output copy to hold a pipeline register if needed

   bh14_w85_9 <= Compressor_3_2_F50_uid49_bh14_uid300_Out0(0);
   bh14_w86_9 <= Compressor_3_2_F50_uid49_bh14_uid300_Out0(1);

   Compressor_23_3_F50_uid41_bh14_uid302_In0 <= "" & bh14_w86_7 & bh14_w86_6 & bh14_w86_5;
   Compressor_23_3_F50_uid41_bh14_uid302_In1 <= "" & bh14_w87_7 & bh14_w87_6;
   Compressor_23_3_F50_uid41_uid302: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid302_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid302_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid302_Out0_copy303);
   Compressor_23_3_F50_uid41_bh14_uid302_Out0 <= Compressor_23_3_F50_uid41_bh14_uid302_Out0_copy303; -- output copy to hold a pipeline register if needed

   bh14_w86_10 <= Compressor_23_3_F50_uid41_bh14_uid302_Out0(0);
   bh14_w87_8 <= Compressor_23_3_F50_uid41_bh14_uid302_Out0(1);
   bh14_w88_8 <= Compressor_23_3_F50_uid41_bh14_uid302_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid304_In0 <= "" & bh14_w88_7 & bh14_w88_6 & bh14_w88_5;
   Compressor_23_3_F50_uid41_bh14_uid304_In1 <= "" & bh14_w89_7 & bh14_w89_6;
   Compressor_23_3_F50_uid41_uid304: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid304_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid304_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid304_Out0_copy305);
   Compressor_23_3_F50_uid41_bh14_uid304_Out0 <= Compressor_23_3_F50_uid41_bh14_uid304_Out0_copy305; -- output copy to hold a pipeline register if needed

   bh14_w88_9 <= Compressor_23_3_F50_uid41_bh14_uid304_Out0(0);
   bh14_w89_8 <= Compressor_23_3_F50_uid41_bh14_uid304_Out0(1);
   bh14_w90_8 <= Compressor_23_3_F50_uid41_bh14_uid304_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid306_In0 <= "" & bh14_w90_7 & bh14_w90_6 & bh14_w90_5;
   Compressor_23_3_F50_uid41_bh14_uid306_In1 <= "" & bh14_w91_7 & bh14_w91_6;
   Compressor_23_3_F50_uid41_uid306: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid306_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid306_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid306_Out0_copy307);
   Compressor_23_3_F50_uid41_bh14_uid306_Out0 <= Compressor_23_3_F50_uid41_bh14_uid306_Out0_copy307; -- output copy to hold a pipeline register if needed

   bh14_w90_9 <= Compressor_23_3_F50_uid41_bh14_uid306_Out0(0);
   bh14_w91_8 <= Compressor_23_3_F50_uid41_bh14_uid306_Out0(1);
   bh14_w92_8 <= Compressor_23_3_F50_uid41_bh14_uid306_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid308_In0 <= "" & bh14_w92_7 & bh14_w92_6 & bh14_w92_5;
   Compressor_23_3_F50_uid41_bh14_uid308_In1 <= "" & bh14_w93_7 & bh14_w93_6;
   Compressor_23_3_F50_uid41_uid308: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid308_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid308_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid308_Out0_copy309);
   Compressor_23_3_F50_uid41_bh14_uid308_Out0 <= Compressor_23_3_F50_uid41_bh14_uid308_Out0_copy309; -- output copy to hold a pipeline register if needed

   bh14_w92_9 <= Compressor_23_3_F50_uid41_bh14_uid308_Out0(0);
   bh14_w93_8 <= Compressor_23_3_F50_uid41_bh14_uid308_Out0(1);
   bh14_w94_7 <= Compressor_23_3_F50_uid41_bh14_uid308_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid310_In0 <= "" & bh14_w94_6 & bh14_w94_5 & bh14_w94_4;
   Compressor_23_3_F50_uid41_bh14_uid310_In1 <= "" & "0" & "0";
   Compressor_23_3_F50_uid41_uid310: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid310_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid310_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid310_Out0_copy311);
   Compressor_23_3_F50_uid41_bh14_uid310_Out0 <= Compressor_23_3_F50_uid41_bh14_uid310_Out0_copy311; -- output copy to hold a pipeline register if needed

   bh14_w94_8 <= Compressor_23_3_F50_uid41_bh14_uid310_Out0(0);
   bh14_w95_7 <= Compressor_23_3_F50_uid41_bh14_uid310_Out0(1);
   bh14_w96_6 <= Compressor_23_3_F50_uid41_bh14_uid310_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid312_In0 <= "" & bh14_w95_6 & bh14_w95_5 & bh14_w95_4;
   Compressor_23_3_F50_uid41_bh14_uid312_In1 <= "" & bh14_w96_5 & bh14_w96_4;
   Compressor_23_3_F50_uid41_uid312: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid312_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid312_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid312_Out0_copy313);
   Compressor_23_3_F50_uid41_bh14_uid312_Out0 <= Compressor_23_3_F50_uid41_bh14_uid312_Out0_copy313; -- output copy to hold a pipeline register if needed

   bh14_w95_8 <= Compressor_23_3_F50_uid41_bh14_uid312_Out0(0);
   bh14_w96_7 <= Compressor_23_3_F50_uid41_bh14_uid312_Out0(1);
   bh14_w97_7 <= Compressor_23_3_F50_uid41_bh14_uid312_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid314_In0 <= "" & bh14_w97_6 & bh14_w97_5 & bh14_w97_4;
   Compressor_23_3_F50_uid41_bh14_uid314_In1 <= "" & bh14_w98_5 & bh14_w98_4;
   Compressor_23_3_F50_uid41_uid314: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid314_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid314_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid314_Out0_copy315);
   Compressor_23_3_F50_uid41_bh14_uid314_Out0 <= Compressor_23_3_F50_uid41_bh14_uid314_Out0_copy315; -- output copy to hold a pipeline register if needed

   bh14_w97_8 <= Compressor_23_3_F50_uid41_bh14_uid314_Out0(0);
   bh14_w98_6 <= Compressor_23_3_F50_uid41_bh14_uid314_Out0(1);
   bh14_w99_7 <= Compressor_23_3_F50_uid41_bh14_uid314_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid316_In0 <= "" & bh14_w99_6 & bh14_w99_5 & bh14_w99_4;
   Compressor_23_3_F50_uid41_bh14_uid316_In1 <= "" & bh14_w100_5 & bh14_w100_4;
   Compressor_23_3_F50_uid41_uid316: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid316_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid316_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid316_Out0_copy317);
   Compressor_23_3_F50_uid41_bh14_uid316_Out0 <= Compressor_23_3_F50_uid41_bh14_uid316_Out0_copy317; -- output copy to hold a pipeline register if needed

   bh14_w99_8 <= Compressor_23_3_F50_uid41_bh14_uid316_Out0(0);
   bh14_w100_6 <= Compressor_23_3_F50_uid41_bh14_uid316_Out0(1);
   bh14_w101_7 <= Compressor_23_3_F50_uid41_bh14_uid316_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid318_In0 <= "" & bh14_w101_6 & bh14_w101_5 & bh14_w101_4;
   Compressor_23_3_F50_uid41_bh14_uid318_In1 <= "" & bh14_w102_5 & bh14_w102_4;
   Compressor_23_3_F50_uid41_uid318: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid318_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid318_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid318_Out0_copy319);
   Compressor_23_3_F50_uid41_bh14_uid318_Out0 <= Compressor_23_3_F50_uid41_bh14_uid318_Out0_copy319; -- output copy to hold a pipeline register if needed

   bh14_w101_8 <= Compressor_23_3_F50_uid41_bh14_uid318_Out0(0);
   bh14_w102_6 <= Compressor_23_3_F50_uid41_bh14_uid318_Out0(1);
   bh14_w103_7 <= Compressor_23_3_F50_uid41_bh14_uid318_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid320_In0 <= "" & bh14_w103_6 & bh14_w103_5 & bh14_w103_4;
   Compressor_23_3_F50_uid41_bh14_uid320_In1 <= "" & bh14_w104_5 & bh14_w104_4;
   Compressor_23_3_F50_uid41_uid320: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid320_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid320_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid320_Out0_copy321);
   Compressor_23_3_F50_uid41_bh14_uid320_Out0 <= Compressor_23_3_F50_uid41_bh14_uid320_Out0_copy321; -- output copy to hold a pipeline register if needed

   bh14_w103_8 <= Compressor_23_3_F50_uid41_bh14_uid320_Out0(0);
   bh14_w104_6 <= Compressor_23_3_F50_uid41_bh14_uid320_Out0(1);
   bh14_w105_7 <= Compressor_23_3_F50_uid41_bh14_uid320_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid322_In0 <= "" & bh14_w105_6 & bh14_w105_5 & bh14_w105_4;
   Compressor_23_3_F50_uid41_bh14_uid322_In1 <= "" & bh14_w106_5 & bh14_w106_4;
   Compressor_23_3_F50_uid41_uid322: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid322_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid322_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid322_Out0_copy323);
   Compressor_23_3_F50_uid41_bh14_uid322_Out0 <= Compressor_23_3_F50_uid41_bh14_uid322_Out0_copy323; -- output copy to hold a pipeline register if needed

   bh14_w105_8 <= Compressor_23_3_F50_uid41_bh14_uid322_Out0(0);
   bh14_w106_6 <= Compressor_23_3_F50_uid41_bh14_uid322_Out0(1);
   bh14_w107_7 <= Compressor_23_3_F50_uid41_bh14_uid322_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid324_In0 <= "" & bh14_w107_6 & bh14_w107_5 & bh14_w107_4;
   Compressor_23_3_F50_uid41_bh14_uid324_In1 <= "" & bh14_w108_3 & bh14_w108_4;
   Compressor_23_3_F50_uid41_uid324: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid324_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid324_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid324_Out0_copy325);
   Compressor_23_3_F50_uid41_bh14_uid324_Out0 <= Compressor_23_3_F50_uid41_bh14_uid324_Out0_copy325; -- output copy to hold a pipeline register if needed

   bh14_w107_8 <= Compressor_23_3_F50_uid41_bh14_uid324_Out0(0);
   bh14_w108_5 <= Compressor_23_3_F50_uid41_bh14_uid324_Out0(1);
   bh14_w109_6 <= Compressor_23_3_F50_uid41_bh14_uid324_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid326_In0 <= "" & bh14_w109_3 & bh14_w109_5 & bh14_w109_4;
   Compressor_23_3_F50_uid41_bh14_uid326_In1 <= "" & bh14_w110_3 & bh14_w110_2;
   Compressor_23_3_F50_uid41_uid326: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid326_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid326_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid326_Out0_copy327);
   Compressor_23_3_F50_uid41_bh14_uid326_Out0 <= Compressor_23_3_F50_uid41_bh14_uid326_Out0_copy327; -- output copy to hold a pipeline register if needed

   bh14_w109_7 <= Compressor_23_3_F50_uid41_bh14_uid326_Out0(0);
   bh14_w110_4 <= Compressor_23_3_F50_uid41_bh14_uid326_Out0(1);
   bh14_w111_4 <= Compressor_23_3_F50_uid41_bh14_uid326_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid328_In0 <= "" & bh14_w111_3 & bh14_w111_2 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid328_In1 <= "" & bh14_w112_2;
   Compressor_14_3_F50_uid63_uid328: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid328_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid328_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid328_Out0_copy329);
   Compressor_14_3_F50_uid63_bh14_uid328_Out0 <= Compressor_14_3_F50_uid63_bh14_uid328_Out0_copy329; -- output copy to hold a pipeline register if needed

   bh14_w111_5 <= Compressor_14_3_F50_uid63_bh14_uid328_Out0(0);
   bh14_w112_3 <= Compressor_14_3_F50_uid63_bh14_uid328_Out0(1);
   bh14_w113_4 <= Compressor_14_3_F50_uid63_bh14_uid328_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid330_In0 <= "" & bh14_w113_3 & bh14_w113_2 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid330_In1 <= "" & bh14_w114_2;
   Compressor_14_3_F50_uid63_uid330: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid330_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid330_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid330_Out0_copy331);
   Compressor_14_3_F50_uid63_bh14_uid330_Out0 <= Compressor_14_3_F50_uid63_bh14_uid330_Out0_copy331; -- output copy to hold a pipeline register if needed

   bh14_w113_5 <= Compressor_14_3_F50_uid63_bh14_uid330_Out0(0);
   bh14_w114_3 <= Compressor_14_3_F50_uid63_bh14_uid330_Out0(1);
   bh14_w115_4 <= Compressor_14_3_F50_uid63_bh14_uid330_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid332_In0 <= "" & bh14_w115_3 & bh14_w115_2 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid332_In1 <= "" & bh14_w116_2;
   Compressor_14_3_F50_uid63_uid332: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid332_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid332_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid332_Out0_copy333);
   Compressor_14_3_F50_uid63_bh14_uid332_Out0 <= Compressor_14_3_F50_uid63_bh14_uid332_Out0_copy333; -- output copy to hold a pipeline register if needed

   bh14_w115_5 <= Compressor_14_3_F50_uid63_bh14_uid332_Out0(0);
   bh14_w116_3 <= Compressor_14_3_F50_uid63_bh14_uid332_Out0(1);
   bh14_w117_4 <= Compressor_14_3_F50_uid63_bh14_uid332_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid334_In0 <= "" & bh14_w117_3 & bh14_w117_2 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid334_In1 <= "" & bh14_w118_2;
   Compressor_14_3_F50_uid63_uid334: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid334_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid334_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid334_Out0_copy335);
   Compressor_14_3_F50_uid63_bh14_uid334_Out0 <= Compressor_14_3_F50_uid63_bh14_uid334_Out0_copy335; -- output copy to hold a pipeline register if needed

   bh14_w117_5 <= Compressor_14_3_F50_uid63_bh14_uid334_Out0(0);
   bh14_w118_3 <= Compressor_14_3_F50_uid63_bh14_uid334_Out0(1);
   bh14_w119_4 <= Compressor_14_3_F50_uid63_bh14_uid334_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid336_In0 <= "" & bh14_w119_3 & bh14_w119_2 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid336_In1 <= "" & bh14_w120_2;
   Compressor_14_3_F50_uid63_uid336: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid336_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid336_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid336_Out0_copy337);
   Compressor_14_3_F50_uid63_bh14_uid336_Out0 <= Compressor_14_3_F50_uid63_bh14_uid336_Out0_copy337; -- output copy to hold a pipeline register if needed

   bh14_w119_5 <= Compressor_14_3_F50_uid63_bh14_uid336_Out0(0);
   bh14_w120_3 <= Compressor_14_3_F50_uid63_bh14_uid336_Out0(1);
   bh14_w121_2 <= Compressor_14_3_F50_uid63_bh14_uid336_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid338_In0 <= "" & bh14_w121_1 & bh14_w121_0 & "0";
   Compressor_3_2_F50_uid49_uid338: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid338_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid338_Out0_copy339);
   Compressor_3_2_F50_uid49_bh14_uid338_Out0 <= Compressor_3_2_F50_uid49_bh14_uid338_Out0_copy339; -- output copy to hold a pipeline register if needed

   bh14_w121_3 <= Compressor_3_2_F50_uid49_bh14_uid338_Out0(0);

   Compressor_14_3_F50_uid63_bh14_uid340_In0 <= "" & bh14_w21_5 & bh14_w21_4 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid340_In1 <= "" & bh14_w22_3;
   Compressor_14_3_F50_uid63_uid340: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid340_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid340_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid340_Out0_copy341);
   Compressor_14_3_F50_uid63_bh14_uid340_Out0 <= Compressor_14_3_F50_uid63_bh14_uid340_Out0_copy341; -- output copy to hold a pipeline register if needed

   bh14_w21_6 <= Compressor_14_3_F50_uid63_bh14_uid340_Out0(0);
   bh14_w22_4 <= Compressor_14_3_F50_uid63_bh14_uid340_Out0(1);
   bh14_w23_6 <= Compressor_14_3_F50_uid63_bh14_uid340_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid342_In0 <= "" & bh14_w23_5 & bh14_w23_4 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid342_In1 <= "" & bh14_w24_5;
   Compressor_14_3_F50_uid63_uid342: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid342_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid342_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid342_Out0_copy343);
   Compressor_14_3_F50_uid63_bh14_uid342_Out0 <= Compressor_14_3_F50_uid63_bh14_uid342_Out0_copy343; -- output copy to hold a pipeline register if needed

   bh14_w23_7 <= Compressor_14_3_F50_uid63_bh14_uid342_Out0(0);
   bh14_w24_6 <= Compressor_14_3_F50_uid63_bh14_uid342_Out0(1);
   bh14_w25_6 <= Compressor_14_3_F50_uid63_bh14_uid342_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid344_In0 <= "" & bh14_w25_5 & bh14_w25_4 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid344_In1 <= "" & bh14_w26_5;
   Compressor_14_3_F50_uid63_uid344: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid344_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid344_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid344_Out0_copy345);
   Compressor_14_3_F50_uid63_bh14_uid344_Out0 <= Compressor_14_3_F50_uid63_bh14_uid344_Out0_copy345; -- output copy to hold a pipeline register if needed

   bh14_w25_7 <= Compressor_14_3_F50_uid63_bh14_uid344_Out0(0);
   bh14_w26_6 <= Compressor_14_3_F50_uid63_bh14_uid344_Out0(1);
   bh14_w27_6 <= Compressor_14_3_F50_uid63_bh14_uid344_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid346_In0 <= "" & bh14_w27_5 & bh14_w27_4 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid346_In1 <= "" & bh14_w28_5;
   Compressor_14_3_F50_uid63_uid346: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid346_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid346_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid346_Out0_copy347);
   Compressor_14_3_F50_uid63_bh14_uid346_Out0 <= Compressor_14_3_F50_uid63_bh14_uid346_Out0_copy347; -- output copy to hold a pipeline register if needed

   bh14_w27_7 <= Compressor_14_3_F50_uid63_bh14_uid346_Out0(0);
   bh14_w28_6 <= Compressor_14_3_F50_uid63_bh14_uid346_Out0(1);
   bh14_w29_6 <= Compressor_14_3_F50_uid63_bh14_uid346_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid348_In0 <= "" & bh14_w29_5 & bh14_w29_4 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid348_In1 <= "" & bh14_w30_5;
   Compressor_14_3_F50_uid63_uid348: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid348_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid348_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid348_Out0_copy349);
   Compressor_14_3_F50_uid63_bh14_uid348_Out0 <= Compressor_14_3_F50_uid63_bh14_uid348_Out0_copy349; -- output copy to hold a pipeline register if needed

   bh14_w29_7 <= Compressor_14_3_F50_uid63_bh14_uid348_Out0(0);
   bh14_w30_6 <= Compressor_14_3_F50_uid63_bh14_uid348_Out0(1);
   bh14_w31_6 <= Compressor_14_3_F50_uid63_bh14_uid348_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid350_In0 <= "" & bh14_w31_5 & bh14_w31_4 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid350_In1 <= "" & bh14_w32_5;
   Compressor_14_3_F50_uid63_uid350: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid350_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid350_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid350_Out0_copy351);
   Compressor_14_3_F50_uid63_bh14_uid350_Out0 <= Compressor_14_3_F50_uid63_bh14_uid350_Out0_copy351; -- output copy to hold a pipeline register if needed

   bh14_w31_7 <= Compressor_14_3_F50_uid63_bh14_uid350_Out0(0);
   bh14_w32_6 <= Compressor_14_3_F50_uid63_bh14_uid350_Out0(1);
   bh14_w33_6 <= Compressor_14_3_F50_uid63_bh14_uid350_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid352_In0 <= "" & bh14_w33_5 & bh14_w33_4 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid352_In1 <= "" & bh14_w34_6;
   Compressor_14_3_F50_uid63_uid352: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid352_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid352_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid352_Out0_copy353);
   Compressor_14_3_F50_uid63_bh14_uid352_Out0 <= Compressor_14_3_F50_uid63_bh14_uid352_Out0_copy353; -- output copy to hold a pipeline register if needed

   bh14_w33_7 <= Compressor_14_3_F50_uid63_bh14_uid352_Out0(0);
   bh14_w34_7 <= Compressor_14_3_F50_uid63_bh14_uid352_Out0(1);
   bh14_w35_8 <= Compressor_14_3_F50_uid63_bh14_uid352_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid354_In0 <= "" & bh14_w35_7 & bh14_w35_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid354_In1 <= "" & bh14_w36_8 & bh14_w36_7;
   Compressor_23_3_F50_uid41_uid354: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid354_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid354_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid354_Out0_copy355);
   Compressor_23_3_F50_uid41_bh14_uid354_Out0 <= Compressor_23_3_F50_uid41_bh14_uid354_Out0_copy355; -- output copy to hold a pipeline register if needed

   bh14_w35_9 <= Compressor_23_3_F50_uid41_bh14_uid354_Out0(0);
   bh14_w36_9 <= Compressor_23_3_F50_uid41_bh14_uid354_Out0(1);
   bh14_w37_7 <= Compressor_23_3_F50_uid41_bh14_uid354_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid356_In0 <= "" & bh14_w38_8 & bh14_w38_7 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid356_In1 <= "" & bh14_w39_6;
   Compressor_14_3_F50_uid63_uid356: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid356_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid356_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid356_Out0_copy357);
   Compressor_14_3_F50_uid63_bh14_uid356_Out0 <= Compressor_14_3_F50_uid63_bh14_uid356_Out0_copy357; -- output copy to hold a pipeline register if needed

   bh14_w38_9 <= Compressor_14_3_F50_uid63_bh14_uid356_Out0(0);
   bh14_w39_7 <= Compressor_14_3_F50_uid63_bh14_uid356_Out0(1);
   bh14_w40_9 <= Compressor_14_3_F50_uid63_bh14_uid356_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid358_In0 <= "" & bh14_w40_8 & bh14_w40_7 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid358_In1 <= "" & bh14_w41_6;
   Compressor_14_3_F50_uid63_uid358: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid358_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid358_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid358_Out0_copy359);
   Compressor_14_3_F50_uid63_bh14_uid358_Out0 <= Compressor_14_3_F50_uid63_bh14_uid358_Out0_copy359; -- output copy to hold a pipeline register if needed

   bh14_w40_10 <= Compressor_14_3_F50_uid63_bh14_uid358_Out0(0);
   bh14_w41_7 <= Compressor_14_3_F50_uid63_bh14_uid358_Out0(1);
   bh14_w42_9 <= Compressor_14_3_F50_uid63_bh14_uid358_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid360_In0 <= "" & bh14_w42_8 & bh14_w42_7 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid360_In1 <= "" & bh14_w43_6;
   Compressor_14_3_F50_uid63_uid360: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid360_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid360_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid360_Out0_copy361);
   Compressor_14_3_F50_uid63_bh14_uid360_Out0 <= Compressor_14_3_F50_uid63_bh14_uid360_Out0_copy361; -- output copy to hold a pipeline register if needed

   bh14_w42_10 <= Compressor_14_3_F50_uid63_bh14_uid360_Out0(0);
   bh14_w43_7 <= Compressor_14_3_F50_uid63_bh14_uid360_Out0(1);
   bh14_w44_9 <= Compressor_14_3_F50_uid63_bh14_uid360_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid362_In0 <= "" & bh14_w44_8 & bh14_w44_7 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid362_In1 <= "" & bh14_w45_6;
   Compressor_14_3_F50_uid63_uid362: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid362_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid362_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid362_Out0_copy363);
   Compressor_14_3_F50_uid63_bh14_uid362_Out0 <= Compressor_14_3_F50_uid63_bh14_uid362_Out0_copy363; -- output copy to hold a pipeline register if needed

   bh14_w44_10 <= Compressor_14_3_F50_uid63_bh14_uid362_Out0(0);
   bh14_w45_7 <= Compressor_14_3_F50_uid63_bh14_uid362_Out0(1);
   bh14_w46_9 <= Compressor_14_3_F50_uid63_bh14_uid362_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid364_In0 <= "" & bh14_w46_8 & bh14_w46_7 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid364_In1 <= "" & bh14_w47_6;
   Compressor_14_3_F50_uid63_uid364: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid364_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid364_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid364_Out0_copy365);
   Compressor_14_3_F50_uid63_bh14_uid364_Out0 <= Compressor_14_3_F50_uid63_bh14_uid364_Out0_copy365; -- output copy to hold a pipeline register if needed

   bh14_w46_10 <= Compressor_14_3_F50_uid63_bh14_uid364_Out0(0);
   bh14_w47_7 <= Compressor_14_3_F50_uid63_bh14_uid364_Out0(1);
   bh14_w48_10 <= Compressor_14_3_F50_uid63_bh14_uid364_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid366_In0 <= "" & bh14_w48_9 & bh14_w48_8 & "0";
   Compressor_23_3_F50_uid41_bh14_uid366_In1 <= "" & bh14_w49_7 & bh14_w49_5;
   Compressor_23_3_F50_uid41_uid366: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid366_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid366_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid366_Out0_copy367);
   Compressor_23_3_F50_uid41_bh14_uid366_Out0 <= Compressor_23_3_F50_uid41_bh14_uid366_Out0_copy367; -- output copy to hold a pipeline register if needed

   bh14_w48_11 <= Compressor_23_3_F50_uid41_bh14_uid366_Out0(0);
   bh14_w49_8 <= Compressor_23_3_F50_uid41_bh14_uid366_Out0(1);
   bh14_w50_10 <= Compressor_23_3_F50_uid41_bh14_uid366_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid368_In0 <= "" & bh14_w50_9 & bh14_w50_8 & "0";
   Compressor_23_3_F50_uid41_bh14_uid368_In1 <= "" & bh14_w51_9 & bh14_w51_10;
   Compressor_23_3_F50_uid41_uid368: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid368_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid368_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid368_Out0_copy369);
   Compressor_23_3_F50_uid41_bh14_uid368_Out0 <= Compressor_23_3_F50_uid41_bh14_uid368_Out0_copy369; -- output copy to hold a pipeline register if needed

   bh14_w50_11 <= Compressor_23_3_F50_uid41_bh14_uid368_Out0(0);
   bh14_w51_11 <= Compressor_23_3_F50_uid41_bh14_uid368_Out0(1);
   bh14_w52_10 <= Compressor_23_3_F50_uid41_bh14_uid368_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid370_In0 <= "" & bh14_w52_8 & bh14_w52_9 & "0";
   Compressor_23_3_F50_uid41_bh14_uid370_In1 <= "" & bh14_w53_10 & bh14_w53_9;
   Compressor_23_3_F50_uid41_uid370: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid370_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid370_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid370_Out0_copy371);
   Compressor_23_3_F50_uid41_bh14_uid370_Out0 <= Compressor_23_3_F50_uid41_bh14_uid370_Out0_copy371; -- output copy to hold a pipeline register if needed

   bh14_w52_11 <= Compressor_23_3_F50_uid41_bh14_uid370_Out0(0);
   bh14_w53_11 <= Compressor_23_3_F50_uid41_bh14_uid370_Out0(1);
   bh14_w54_10 <= Compressor_23_3_F50_uid41_bh14_uid370_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid372_In0 <= "" & bh14_w54_9 & bh14_w54_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid372_In1 <= "" & bh14_w55_10 & bh14_w55_9;
   Compressor_23_3_F50_uid41_uid372: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid372_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid372_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid372_Out0_copy373);
   Compressor_23_3_F50_uid41_bh14_uid372_Out0 <= Compressor_23_3_F50_uid41_bh14_uid372_Out0_copy373; -- output copy to hold a pipeline register if needed

   bh14_w54_11 <= Compressor_23_3_F50_uid41_bh14_uid372_Out0(0);
   bh14_w55_11 <= Compressor_23_3_F50_uid41_bh14_uid372_Out0(1);
   bh14_w56_10 <= Compressor_23_3_F50_uid41_bh14_uid372_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid374_In0 <= "" & bh14_w56_9 & bh14_w56_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid374_In1 <= "" & bh14_w57_10 & bh14_w57_9;
   Compressor_23_3_F50_uid41_uid374: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid374_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid374_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid374_Out0_copy375);
   Compressor_23_3_F50_uid41_bh14_uid374_Out0 <= Compressor_23_3_F50_uid41_bh14_uid374_Out0_copy375; -- output copy to hold a pipeline register if needed

   bh14_w56_11 <= Compressor_23_3_F50_uid41_bh14_uid374_Out0(0);
   bh14_w57_11 <= Compressor_23_3_F50_uid41_bh14_uid374_Out0(1);
   bh14_w58_10 <= Compressor_23_3_F50_uid41_bh14_uid374_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid376_In0 <= "" & bh14_w58_9 & bh14_w58_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid376_In1 <= "" & bh14_w59_10 & bh14_w59_9;
   Compressor_23_3_F50_uid41_uid376: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid376_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid376_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid376_Out0_copy377);
   Compressor_23_3_F50_uid41_bh14_uid376_Out0 <= Compressor_23_3_F50_uid41_bh14_uid376_Out0_copy377; -- output copy to hold a pipeline register if needed

   bh14_w58_11 <= Compressor_23_3_F50_uid41_bh14_uid376_Out0(0);
   bh14_w59_11 <= Compressor_23_3_F50_uid41_bh14_uid376_Out0(1);
   bh14_w60_10 <= Compressor_23_3_F50_uid41_bh14_uid376_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid378_In0 <= "" & bh14_w60_9 & bh14_w60_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid378_In1 <= "" & bh14_w61_10 & bh14_w61_9;
   Compressor_23_3_F50_uid41_uid378: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid378_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid378_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid378_Out0_copy379);
   Compressor_23_3_F50_uid41_bh14_uid378_Out0 <= Compressor_23_3_F50_uid41_bh14_uid378_Out0_copy379; -- output copy to hold a pipeline register if needed

   bh14_w60_11 <= Compressor_23_3_F50_uid41_bh14_uid378_Out0(0);
   bh14_w61_11 <= Compressor_23_3_F50_uid41_bh14_uid378_Out0(1);
   bh14_w62_10 <= Compressor_23_3_F50_uid41_bh14_uid378_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid380_In0 <= "" & bh14_w62_9 & bh14_w62_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid380_In1 <= "" & bh14_w63_10 & bh14_w63_9;
   Compressor_23_3_F50_uid41_uid380: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid380_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid380_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid380_Out0_copy381);
   Compressor_23_3_F50_uid41_bh14_uid380_Out0 <= Compressor_23_3_F50_uid41_bh14_uid380_Out0_copy381; -- output copy to hold a pipeline register if needed

   bh14_w62_11 <= Compressor_23_3_F50_uid41_bh14_uid380_Out0(0);
   bh14_w63_11 <= Compressor_23_3_F50_uid41_bh14_uid380_Out0(1);
   bh14_w64_10 <= Compressor_23_3_F50_uid41_bh14_uid380_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid382_In0 <= "" & bh14_w64_9 & bh14_w64_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid382_In1 <= "" & bh14_w65_10 & bh14_w65_9;
   Compressor_23_3_F50_uid41_uid382: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid382_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid382_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid382_Out0_copy383);
   Compressor_23_3_F50_uid41_bh14_uid382_Out0 <= Compressor_23_3_F50_uid41_bh14_uid382_Out0_copy383; -- output copy to hold a pipeline register if needed

   bh14_w64_11 <= Compressor_23_3_F50_uid41_bh14_uid382_Out0(0);
   bh14_w65_11 <= Compressor_23_3_F50_uid41_bh14_uid382_Out0(1);
   bh14_w66_10 <= Compressor_23_3_F50_uid41_bh14_uid382_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid384_In0 <= "" & bh14_w66_9 & bh14_w66_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid384_In1 <= "" & bh14_w67_10 & bh14_w67_9;
   Compressor_23_3_F50_uid41_uid384: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid384_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid384_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid384_Out0_copy385);
   Compressor_23_3_F50_uid41_bh14_uid384_Out0 <= Compressor_23_3_F50_uid41_bh14_uid384_Out0_copy385; -- output copy to hold a pipeline register if needed

   bh14_w66_11 <= Compressor_23_3_F50_uid41_bh14_uid384_Out0(0);
   bh14_w67_11 <= Compressor_23_3_F50_uid41_bh14_uid384_Out0(1);
   bh14_w68_10 <= Compressor_23_3_F50_uid41_bh14_uid384_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid386_In0 <= "" & bh14_w68_9 & bh14_w68_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid386_In1 <= "" & bh14_w69_10 & bh14_w69_9;
   Compressor_23_3_F50_uid41_uid386: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid386_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid386_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid386_Out0_copy387);
   Compressor_23_3_F50_uid41_bh14_uid386_Out0 <= Compressor_23_3_F50_uid41_bh14_uid386_Out0_copy387; -- output copy to hold a pipeline register if needed

   bh14_w68_11 <= Compressor_23_3_F50_uid41_bh14_uid386_Out0(0);
   bh14_w69_11 <= Compressor_23_3_F50_uid41_bh14_uid386_Out0(1);
   bh14_w70_10 <= Compressor_23_3_F50_uid41_bh14_uid386_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid388_In0 <= "" & bh14_w70_9 & bh14_w70_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid388_In1 <= "" & bh14_w71_10 & bh14_w71_9;
   Compressor_23_3_F50_uid41_uid388: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid388_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid388_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid388_Out0_copy389);
   Compressor_23_3_F50_uid41_bh14_uid388_Out0 <= Compressor_23_3_F50_uid41_bh14_uid388_Out0_copy389; -- output copy to hold a pipeline register if needed

   bh14_w70_11 <= Compressor_23_3_F50_uid41_bh14_uid388_Out0(0);
   bh14_w71_11 <= Compressor_23_3_F50_uid41_bh14_uid388_Out0(1);
   bh14_w72_10 <= Compressor_23_3_F50_uid41_bh14_uid388_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid390_In0 <= "" & bh14_w72_9 & bh14_w72_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid390_In1 <= "" & bh14_w73_10 & bh14_w73_9;
   Compressor_23_3_F50_uid41_uid390: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid390_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid390_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid390_Out0_copy391);
   Compressor_23_3_F50_uid41_bh14_uid390_Out0 <= Compressor_23_3_F50_uid41_bh14_uid390_Out0_copy391; -- output copy to hold a pipeline register if needed

   bh14_w72_11 <= Compressor_23_3_F50_uid41_bh14_uid390_Out0(0);
   bh14_w73_11 <= Compressor_23_3_F50_uid41_bh14_uid390_Out0(1);
   bh14_w74_10 <= Compressor_23_3_F50_uid41_bh14_uid390_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid392_In0 <= "" & bh14_w74_9 & bh14_w74_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid392_In1 <= "" & bh14_w75_10 & bh14_w75_9;
   Compressor_23_3_F50_uid41_uid392: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid392_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid392_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid392_Out0_copy393);
   Compressor_23_3_F50_uid41_bh14_uid392_Out0 <= Compressor_23_3_F50_uid41_bh14_uid392_Out0_copy393; -- output copy to hold a pipeline register if needed

   bh14_w74_11 <= Compressor_23_3_F50_uid41_bh14_uid392_Out0(0);
   bh14_w75_11 <= Compressor_23_3_F50_uid41_bh14_uid392_Out0(1);
   bh14_w76_10 <= Compressor_23_3_F50_uid41_bh14_uid392_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid394_In0 <= "" & bh14_w76_9 & bh14_w76_6 & "0";
   Compressor_23_3_F50_uid41_bh14_uid394_In1 <= "" & bh14_w77_11 & bh14_w77_10;
   Compressor_23_3_F50_uid41_uid394: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid394_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid394_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid394_Out0_copy395);
   Compressor_23_3_F50_uid41_bh14_uid394_Out0 <= Compressor_23_3_F50_uid41_bh14_uid394_Out0_copy395; -- output copy to hold a pipeline register if needed

   bh14_w76_11 <= Compressor_23_3_F50_uid41_bh14_uid394_Out0(0);
   bh14_w77_12 <= Compressor_23_3_F50_uid41_bh14_uid394_Out0(1);
   bh14_w78_11 <= Compressor_23_3_F50_uid41_bh14_uid394_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid396_In0 <= "" & bh14_w78_9 & bh14_w78_10 & "0";
   Compressor_3_2_F50_uid49_uid396: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid396_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid396_Out0_copy397);
   Compressor_3_2_F50_uid49_bh14_uid396_Out0 <= Compressor_3_2_F50_uid49_bh14_uid396_Out0_copy397; -- output copy to hold a pipeline register if needed

   bh14_w78_12 <= Compressor_3_2_F50_uid49_bh14_uid396_Out0(0);
   bh14_w79_12 <= Compressor_3_2_F50_uid49_bh14_uid396_Out0(1);

   Compressor_23_3_F50_uid41_bh14_uid398_In0 <= "" & bh14_w79_9 & bh14_w79_11 & bh14_w79_10;
   Compressor_23_3_F50_uid41_bh14_uid398_In1 <= "" & bh14_w80_9 & bh14_w80_6;
   Compressor_23_3_F50_uid41_uid398: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid398_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid398_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid398_Out0_copy399);
   Compressor_23_3_F50_uid41_bh14_uid398_Out0 <= Compressor_23_3_F50_uid41_bh14_uid398_Out0_copy399; -- output copy to hold a pipeline register if needed

   bh14_w79_13 <= Compressor_23_3_F50_uid41_bh14_uid398_Out0(0);
   bh14_w80_10 <= Compressor_23_3_F50_uid41_bh14_uid398_Out0(1);
   bh14_w81_11 <= Compressor_23_3_F50_uid41_bh14_uid398_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid400_In0 <= "" & bh14_w81_10 & bh14_w81_9 & "0";
   Compressor_23_3_F50_uid41_bh14_uid400_In1 <= "" & bh14_w82_9 & bh14_w82_6;
   Compressor_23_3_F50_uid41_uid400: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid400_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid400_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid400_Out0_copy401);
   Compressor_23_3_F50_uid41_bh14_uid400_Out0 <= Compressor_23_3_F50_uid41_bh14_uid400_Out0_copy401; -- output copy to hold a pipeline register if needed

   bh14_w81_12 <= Compressor_23_3_F50_uid41_bh14_uid400_Out0(0);
   bh14_w82_10 <= Compressor_23_3_F50_uid41_bh14_uid400_Out0(1);
   bh14_w83_11 <= Compressor_23_3_F50_uid41_bh14_uid400_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid402_In0 <= "" & bh14_w83_10 & bh14_w83_9 & "0";
   Compressor_23_3_F50_uid41_bh14_uid402_In1 <= "" & bh14_w84_9 & bh14_w84_8;
   Compressor_23_3_F50_uid41_uid402: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid402_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid402_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid402_Out0_copy403);
   Compressor_23_3_F50_uid41_bh14_uid402_Out0 <= Compressor_23_3_F50_uid41_bh14_uid402_Out0_copy403; -- output copy to hold a pipeline register if needed

   bh14_w83_12 <= Compressor_23_3_F50_uid41_bh14_uid402_Out0(0);
   bh14_w84_10 <= Compressor_23_3_F50_uid41_bh14_uid402_Out0(1);
   bh14_w85_10 <= Compressor_23_3_F50_uid41_bh14_uid402_Out0(2);

   Compressor_3_2_F50_uid49_bh14_uid404_In0 <= "" & bh14_w85_8 & bh14_w85_9 & "0";
   Compressor_3_2_F50_uid49_uid404: Compressor_3_2_F50_uid49
      port map ( X0 => Compressor_3_2_F50_uid49_bh14_uid404_In0,
                 R => Compressor_3_2_F50_uid49_bh14_uid404_Out0_copy405);
   Compressor_3_2_F50_uid49_bh14_uid404_Out0 <= Compressor_3_2_F50_uid49_bh14_uid404_Out0_copy405; -- output copy to hold a pipeline register if needed

   bh14_w85_11 <= Compressor_3_2_F50_uid49_bh14_uid404_Out0(0);
   bh14_w86_11 <= Compressor_3_2_F50_uid49_bh14_uid404_Out0(1);

   Compressor_23_3_F50_uid41_bh14_uid406_In0 <= "" & bh14_w86_8 & bh14_w86_10 & bh14_w86_9;
   Compressor_23_3_F50_uid41_bh14_uid406_In1 <= "" & bh14_w87_8 & bh14_w87_5;
   Compressor_23_3_F50_uid41_uid406: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid406_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid406_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid406_Out0_copy407);
   Compressor_23_3_F50_uid41_bh14_uid406_Out0 <= Compressor_23_3_F50_uid41_bh14_uid406_Out0_copy407; -- output copy to hold a pipeline register if needed

   bh14_w86_12 <= Compressor_23_3_F50_uid41_bh14_uid406_Out0(0);
   bh14_w87_9 <= Compressor_23_3_F50_uid41_bh14_uid406_Out0(1);
   bh14_w88_10 <= Compressor_23_3_F50_uid41_bh14_uid406_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid408_In0 <= "" & bh14_w88_9 & bh14_w88_8 & "0";
   Compressor_23_3_F50_uid41_bh14_uid408_In1 <= "" & bh14_w89_8 & bh14_w89_5;
   Compressor_23_3_F50_uid41_uid408: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid408_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid408_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid408_Out0_copy409);
   Compressor_23_3_F50_uid41_bh14_uid408_Out0 <= Compressor_23_3_F50_uid41_bh14_uid408_Out0_copy409; -- output copy to hold a pipeline register if needed

   bh14_w88_11 <= Compressor_23_3_F50_uid41_bh14_uid408_Out0(0);
   bh14_w89_9 <= Compressor_23_3_F50_uid41_bh14_uid408_Out0(1);
   bh14_w90_10 <= Compressor_23_3_F50_uid41_bh14_uid408_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid410_In0 <= "" & bh14_w90_9 & bh14_w90_8 & "0";
   Compressor_23_3_F50_uid41_bh14_uid410_In1 <= "" & bh14_w91_8 & bh14_w91_5;
   Compressor_23_3_F50_uid41_uid410: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid410_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid410_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid410_Out0_copy411);
   Compressor_23_3_F50_uid41_bh14_uid410_Out0 <= Compressor_23_3_F50_uid41_bh14_uid410_Out0_copy411; -- output copy to hold a pipeline register if needed

   bh14_w90_11 <= Compressor_23_3_F50_uid41_bh14_uid410_Out0(0);
   bh14_w91_9 <= Compressor_23_3_F50_uid41_bh14_uid410_Out0(1);
   bh14_w92_10 <= Compressor_23_3_F50_uid41_bh14_uid410_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid412_In0 <= "" & bh14_w92_9 & bh14_w92_8 & "0";
   Compressor_23_3_F50_uid41_bh14_uid412_In1 <= "" & bh14_w93_8 & bh14_w93_5;
   Compressor_23_3_F50_uid41_uid412: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid412_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid412_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid412_Out0_copy413);
   Compressor_23_3_F50_uid41_bh14_uid412_Out0 <= Compressor_23_3_F50_uid41_bh14_uid412_Out0_copy413; -- output copy to hold a pipeline register if needed

   bh14_w92_11 <= Compressor_23_3_F50_uid41_bh14_uid412_Out0(0);
   bh14_w93_9 <= Compressor_23_3_F50_uid41_bh14_uid412_Out0(1);
   bh14_w94_9 <= Compressor_23_3_F50_uid41_bh14_uid412_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid414_In0 <= "" & bh14_w94_8 & bh14_w94_7 & "0";
   Compressor_23_3_F50_uid41_bh14_uid414_In1 <= "" & bh14_w95_7 & bh14_w95_8;
   Compressor_23_3_F50_uid41_uid414: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid414_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid414_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid414_Out0_copy415);
   Compressor_23_3_F50_uid41_bh14_uid414_Out0 <= Compressor_23_3_F50_uid41_bh14_uid414_Out0_copy415; -- output copy to hold a pipeline register if needed

   bh14_w94_10 <= Compressor_23_3_F50_uid41_bh14_uid414_Out0(0);
   bh14_w95_9 <= Compressor_23_3_F50_uid41_bh14_uid414_Out0(1);
   bh14_w96_8 <= Compressor_23_3_F50_uid41_bh14_uid414_Out0(2);

   Compressor_23_3_F50_uid41_bh14_uid416_In0 <= "" & bh14_w96_6 & bh14_w96_7 & "0";
   Compressor_23_3_F50_uid41_bh14_uid416_In1 <= "" & bh14_w97_8 & bh14_w97_7;
   Compressor_23_3_F50_uid41_uid416: Compressor_23_3_F50_uid41
      port map ( X0 => Compressor_23_3_F50_uid41_bh14_uid416_In0,
                 X1 => Compressor_23_3_F50_uid41_bh14_uid416_In1,
                 R => Compressor_23_3_F50_uid41_bh14_uid416_Out0_copy417);
   Compressor_23_3_F50_uid41_bh14_uid416_Out0 <= Compressor_23_3_F50_uid41_bh14_uid416_Out0_copy417; -- output copy to hold a pipeline register if needed

   bh14_w96_9 <= Compressor_23_3_F50_uid41_bh14_uid416_Out0(0);
   bh14_w97_9 <= Compressor_23_3_F50_uid41_bh14_uid416_Out0(1);
   bh14_w98_7 <= Compressor_23_3_F50_uid41_bh14_uid416_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid418_In0 <= "" & bh14_w99_8 & bh14_w99_7 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid418_In1 <= "" & bh14_w100_6;
   Compressor_14_3_F50_uid63_uid418: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid418_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid418_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid418_Out0_copy419);
   Compressor_14_3_F50_uid63_bh14_uid418_Out0 <= Compressor_14_3_F50_uid63_bh14_uid418_Out0_copy419; -- output copy to hold a pipeline register if needed

   bh14_w99_9 <= Compressor_14_3_F50_uid63_bh14_uid418_Out0(0);
   bh14_w100_7 <= Compressor_14_3_F50_uid63_bh14_uid418_Out0(1);
   bh14_w101_9 <= Compressor_14_3_F50_uid63_bh14_uid418_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid420_In0 <= "" & bh14_w101_8 & bh14_w101_7 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid420_In1 <= "" & bh14_w102_6;
   Compressor_14_3_F50_uid63_uid420: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid420_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid420_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid420_Out0_copy421);
   Compressor_14_3_F50_uid63_bh14_uid420_Out0 <= Compressor_14_3_F50_uid63_bh14_uid420_Out0_copy421; -- output copy to hold a pipeline register if needed

   bh14_w101_10 <= Compressor_14_3_F50_uid63_bh14_uid420_Out0(0);
   bh14_w102_7 <= Compressor_14_3_F50_uid63_bh14_uid420_Out0(1);
   bh14_w103_9 <= Compressor_14_3_F50_uid63_bh14_uid420_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid422_In0 <= "" & bh14_w103_8 & bh14_w103_7 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid422_In1 <= "" & bh14_w104_6;
   Compressor_14_3_F50_uid63_uid422: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid422_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid422_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid422_Out0_copy423);
   Compressor_14_3_F50_uid63_bh14_uid422_Out0 <= Compressor_14_3_F50_uid63_bh14_uid422_Out0_copy423; -- output copy to hold a pipeline register if needed

   bh14_w103_10 <= Compressor_14_3_F50_uid63_bh14_uid422_Out0(0);
   bh14_w104_7 <= Compressor_14_3_F50_uid63_bh14_uid422_Out0(1);
   bh14_w105_9 <= Compressor_14_3_F50_uid63_bh14_uid422_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid424_In0 <= "" & bh14_w105_8 & bh14_w105_7 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid424_In1 <= "" & bh14_w106_6;
   Compressor_14_3_F50_uid63_uid424: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid424_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid424_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid424_Out0_copy425);
   Compressor_14_3_F50_uid63_bh14_uid424_Out0 <= Compressor_14_3_F50_uid63_bh14_uid424_Out0_copy425; -- output copy to hold a pipeline register if needed

   bh14_w105_10 <= Compressor_14_3_F50_uid63_bh14_uid424_Out0(0);
   bh14_w106_7 <= Compressor_14_3_F50_uid63_bh14_uid424_Out0(1);
   bh14_w107_9 <= Compressor_14_3_F50_uid63_bh14_uid424_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid426_In0 <= "" & bh14_w107_8 & bh14_w107_7 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid426_In1 <= "" & bh14_w108_5;
   Compressor_14_3_F50_uid63_uid426: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid426_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid426_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid426_Out0_copy427);
   Compressor_14_3_F50_uid63_bh14_uid426_Out0 <= Compressor_14_3_F50_uid63_bh14_uid426_Out0_copy427; -- output copy to hold a pipeline register if needed

   bh14_w107_10 <= Compressor_14_3_F50_uid63_bh14_uid426_Out0(0);
   bh14_w108_6 <= Compressor_14_3_F50_uid63_bh14_uid426_Out0(1);
   bh14_w109_8 <= Compressor_14_3_F50_uid63_bh14_uid426_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid428_In0 <= "" & bh14_w109_6 & bh14_w109_7 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid428_In1 <= "" & bh14_w110_4;
   Compressor_14_3_F50_uid63_uid428: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid428_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid428_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid428_Out0_copy429);
   Compressor_14_3_F50_uid63_bh14_uid428_Out0 <= Compressor_14_3_F50_uid63_bh14_uid428_Out0_copy429; -- output copy to hold a pipeline register if needed

   bh14_w109_9 <= Compressor_14_3_F50_uid63_bh14_uid428_Out0(0);
   bh14_w110_5 <= Compressor_14_3_F50_uid63_bh14_uid428_Out0(1);
   bh14_w111_6 <= Compressor_14_3_F50_uid63_bh14_uid428_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid430_In0 <= "" & bh14_w111_4 & bh14_w111_5 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid430_In1 <= "" & bh14_w112_3;
   Compressor_14_3_F50_uid63_uid430: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid430_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid430_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid430_Out0_copy431);
   Compressor_14_3_F50_uid63_bh14_uid430_Out0 <= Compressor_14_3_F50_uid63_bh14_uid430_Out0_copy431; -- output copy to hold a pipeline register if needed

   bh14_w111_7 <= Compressor_14_3_F50_uid63_bh14_uid430_Out0(0);
   bh14_w112_4 <= Compressor_14_3_F50_uid63_bh14_uid430_Out0(1);
   bh14_w113_6 <= Compressor_14_3_F50_uid63_bh14_uid430_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid432_In0 <= "" & bh14_w113_5 & bh14_w113_4 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid432_In1 <= "" & bh14_w114_3;
   Compressor_14_3_F50_uid63_uid432: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid432_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid432_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid432_Out0_copy433);
   Compressor_14_3_F50_uid63_bh14_uid432_Out0 <= Compressor_14_3_F50_uid63_bh14_uid432_Out0_copy433; -- output copy to hold a pipeline register if needed

   bh14_w113_7 <= Compressor_14_3_F50_uid63_bh14_uid432_Out0(0);
   bh14_w114_4 <= Compressor_14_3_F50_uid63_bh14_uid432_Out0(1);
   bh14_w115_6 <= Compressor_14_3_F50_uid63_bh14_uid432_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid434_In0 <= "" & bh14_w115_5 & bh14_w115_4 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid434_In1 <= "" & bh14_w116_3;
   Compressor_14_3_F50_uid63_uid434: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid434_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid434_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid434_Out0_copy435);
   Compressor_14_3_F50_uid63_bh14_uid434_Out0 <= Compressor_14_3_F50_uid63_bh14_uid434_Out0_copy435; -- output copy to hold a pipeline register if needed

   bh14_w115_7 <= Compressor_14_3_F50_uid63_bh14_uid434_Out0(0);
   bh14_w116_4 <= Compressor_14_3_F50_uid63_bh14_uid434_Out0(1);
   bh14_w117_6 <= Compressor_14_3_F50_uid63_bh14_uid434_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid436_In0 <= "" & bh14_w117_5 & bh14_w117_4 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid436_In1 <= "" & bh14_w118_3;
   Compressor_14_3_F50_uid63_uid436: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid436_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid436_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid436_Out0_copy437);
   Compressor_14_3_F50_uid63_bh14_uid436_Out0 <= Compressor_14_3_F50_uid63_bh14_uid436_Out0_copy437; -- output copy to hold a pipeline register if needed

   bh14_w117_7 <= Compressor_14_3_F50_uid63_bh14_uid436_Out0(0);
   bh14_w118_4 <= Compressor_14_3_F50_uid63_bh14_uid436_Out0(1);
   bh14_w119_6 <= Compressor_14_3_F50_uid63_bh14_uid436_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid438_In0 <= "" & bh14_w119_5 & bh14_w119_4 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid438_In1 <= "" & bh14_w120_3;
   Compressor_14_3_F50_uid63_uid438: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid438_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid438_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid438_Out0_copy439);
   Compressor_14_3_F50_uid63_bh14_uid438_Out0 <= Compressor_14_3_F50_uid63_bh14_uid438_Out0_copy439; -- output copy to hold a pipeline register if needed

   bh14_w119_7 <= Compressor_14_3_F50_uid63_bh14_uid438_Out0(0);
   bh14_w120_4 <= Compressor_14_3_F50_uid63_bh14_uid438_Out0(1);
   bh14_w121_4 <= Compressor_14_3_F50_uid63_bh14_uid438_Out0(2);

   Compressor_14_3_F50_uid63_bh14_uid440_In0 <= "" & bh14_w121_3 & bh14_w121_2 & "0" & "0";
   Compressor_14_3_F50_uid63_bh14_uid440_In1 <= "" & "0";
   Compressor_14_3_F50_uid63_uid440: Compressor_14_3_F50_uid63
      port map ( X0 => Compressor_14_3_F50_uid63_bh14_uid440_In0,
                 X1 => Compressor_14_3_F50_uid63_bh14_uid440_In1,
                 R => Compressor_14_3_F50_uid63_bh14_uid440_Out0_copy441);
   Compressor_14_3_F50_uid63_bh14_uid440_Out0 <= Compressor_14_3_F50_uid63_bh14_uid440_Out0_copy441; -- output copy to hold a pipeline register if needed

   bh14_w121_5 <= Compressor_14_3_F50_uid63_bh14_uid440_Out0(0);
   tmp_bitheapResult_bh14_22 <= bh14_w22_4 & bh14_w21_6 & bh14_w20_3 & bh14_w19_4 & bh14_w18_2 & bh14_w17_2 & bh14_w16_0 & bh14_w15_0 & bh14_w14_0 & bh14_w13_0 & bh14_w12_0 & bh14_w11_0 & bh14_w10_0 & bh14_w9_0 & bh14_w8_0 & bh14_w7_0 & bh14_w6_0 & bh14_w5_0 & bh14_w4_0 & bh14_w3_0 & bh14_w2_0 & bh14_w1_0 & bh14_w0_0;

   bitheapFinalAdd_bh14_In0 <= "0" & bh14_w121_5 & bh14_w120_4 & bh14_w119_7 & bh14_w118_4 & bh14_w117_7 & bh14_w116_4 & bh14_w115_7 & bh14_w114_4 & bh14_w113_6 & bh14_w112_4 & bh14_w111_6 & bh14_w110_5 & bh14_w109_8 & bh14_w108_6 & bh14_w107_10 & bh14_w106_7 & bh14_w105_10 & bh14_w104_7 & bh14_w103_10 & bh14_w102_7 & bh14_w101_10 & bh14_w100_7 & bh14_w99_9 & bh14_w98_7 & bh14_w97_9 & bh14_w96_8 & bh14_w95_9 & bh14_w94_10 & bh14_w93_9 & bh14_w92_11 & bh14_w91_9 & bh14_w90_11 & bh14_w89_9 & bh14_w88_10 & bh14_w87_9 & bh14_w86_11 & bh14_w85_10 & bh14_w84_10 & bh14_w83_12 & bh14_w82_10 & bh14_w81_11 & bh14_w80_10 & bh14_w79_12 & bh14_w78_11 & bh14_w77_12 & bh14_w76_11 & bh14_w75_11 & bh14_w74_11 & bh14_w73_11 & bh14_w72_11 & bh14_w71_11 & bh14_w70_11 & bh14_w69_11 & bh14_w68_11 & bh14_w67_11 & bh14_w66_11 & bh14_w65_11 & bh14_w64_11 & bh14_w63_11 & bh14_w62_11 & bh14_w61_11 & bh14_w60_11 & bh14_w59_11 & bh14_w58_11 & bh14_w57_11 & bh14_w56_11 & bh14_w55_11 & bh14_w54_10 & bh14_w53_11 & bh14_w52_10 & bh14_w51_11 & bh14_w50_11 & bh14_w49_8 & bh14_w48_11 & bh14_w47_7 & bh14_w46_10 & bh14_w45_7 & bh14_w44_10 & bh14_w43_7 & bh14_w42_10 & bh14_w41_7 & bh14_w40_10 & bh14_w39_7 & bh14_w38_9 & bh14_w37_7 & bh14_w36_9 & bh14_w35_9 & bh14_w34_7 & bh14_w33_7 & bh14_w32_6 & bh14_w31_7 & bh14_w30_6 & bh14_w29_7 & bh14_w28_6 & bh14_w27_7 & bh14_w26_6 & bh14_w25_7 & bh14_w24_6 & bh14_w23_7;
   bitheapFinalAdd_bh14_In1 <= "0" & bh14_w121_4 & "0" & bh14_w119_6 & "0" & bh14_w117_6 & "0" & bh14_w115_6 & "0" & bh14_w113_7 & "0" & bh14_w111_7 & "0" & bh14_w109_9 & "0" & bh14_w107_9 & "0" & bh14_w105_9 & "0" & bh14_w103_9 & "0" & bh14_w101_9 & "0" & "0" & bh14_w98_6 & "0" & bh14_w96_9 & "0" & bh14_w94_9 & "0" & bh14_w92_10 & "0" & bh14_w90_10 & "0" & bh14_w88_11 & "0" & bh14_w86_12 & bh14_w85_11 & "0" & bh14_w83_11 & "0" & bh14_w81_12 & "0" & bh14_w79_13 & bh14_w78_12 & "0" & bh14_w76_10 & "0" & bh14_w74_10 & "0" & bh14_w72_10 & "0" & bh14_w70_10 & "0" & bh14_w68_10 & "0" & bh14_w66_10 & "0" & bh14_w64_10 & "0" & bh14_w62_10 & "0" & bh14_w60_10 & "0" & bh14_w58_10 & "0" & bh14_w56_10 & "0" & bh14_w54_11 & "0" & bh14_w52_11 & "0" & bh14_w50_10 & "0" & bh14_w48_10 & "0" & bh14_w46_9 & "0" & bh14_w44_9 & "0" & bh14_w42_9 & "0" & bh14_w40_9 & "0" & "0" & bh14_w37_6 & "0" & bh14_w35_8 & "0" & bh14_w33_6 & "0" & bh14_w31_6 & "0" & bh14_w29_6 & "0" & bh14_w27_6 & "0" & bh14_w25_6 & "0" & bh14_w23_6;
   bitheapFinalAdd_bh14_Cin <= '0';

   bitheapFinalAdd_bh14: IntAdder_100_F50_uid443
      port map ( clk  => clk,
                 Cin => bitheapFinalAdd_bh14_Cin,
                 X => bitheapFinalAdd_bh14_In0,
                 Y => bitheapFinalAdd_bh14_In1,
                 R => bitheapFinalAdd_bh14_Out);
   bitheapResult_bh14 <= bitheapFinalAdd_bh14_Out(98 downto 0) & tmp_bitheapResult_bh14_22;
   R <= bitheapResult_bh14(121 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_10_F50_uid445
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_10_F50_uid445 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : in  std_logic_vector(9 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of IntAdder_10_F50_uid445 is
signal Rtmp :  std_logic_vector(9 downto 0);
begin
   Rtmp <= X + Y + Cin;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_10_F50_uid448
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_10_F50_uid448 is
    port (clk : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : in  std_logic_vector(9 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of IntAdder_10_F50_uid448 is
signal Rtmp :  std_logic_vector(9 downto 0);
begin
   Rtmp <= X + Y + Cin;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                           IntAdder_9_F50_uid450
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_9_F50_uid450 is
    port (clk : in std_logic;
          X : in  std_logic_vector(8 downto 0);
          Y : in  std_logic_vector(8 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(8 downto 0)   );
end entity;

architecture arch of IntAdder_9_F50_uid450 is
signal Rtmp :  std_logic_vector(8 downto 0);
begin
   Rtmp <= X + Y + Cin;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                   RightShifter616_by_max_496_F50_uid452
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca (2008-2011), Florent de Dinechin (2008-2019)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X S padBit
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifter616_by_max_496_F50_uid452 is
    port (clk : in std_logic;
          X : in  std_logic_vector(615 downto 0);
          S : in  std_logic_vector(8 downto 0);
          padBit : in  std_logic;
          R : out  std_logic_vector(615 downto 0)   );
end entity;

architecture arch of RightShifter616_by_max_496_F50_uid452 is
signal ps, ps_d1, ps_d2, ps_d3 :  std_logic_vector(8 downto 0);
signal level0 :  std_logic_vector(615 downto 0);
signal level1, level1_d1 :  std_logic_vector(616 downto 0);
signal level2 :  std_logic_vector(618 downto 0);
signal level3 :  std_logic_vector(622 downto 0);
signal level4 :  std_logic_vector(630 downto 0);
signal level5, level5_d1 :  std_logic_vector(646 downto 0);
signal level6 :  std_logic_vector(678 downto 0);
signal level7, level7_d1 :  std_logic_vector(742 downto 0);
signal level8 :  std_logic_vector(870 downto 0);
signal level9 :  std_logic_vector(1126 downto 0);
signal padBit_d1, padBit_d2, padBit_d3 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            ps_d2 <=  ps_d1;
            ps_d3 <=  ps_d2;
            level1_d1 <=  level1;
            level5_d1 <=  level5;
            level7_d1 <=  level7;
            padBit_d1 <=  padBit;
            padBit_d2 <=  padBit_d1;
            padBit_d3 <=  padBit_d2;
         end if;
      end process;
   ps<= S;
   level0<= X;
   level1 <=  (0 downto 0 => padBit) & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2 <=  (1 downto 0 => padBit_d1) & level1_d1 when ps_d1(1) = '1' else    level1_d1 & (1 downto 0 => '0');
   level3 <=  (3 downto 0 => padBit_d1) & level2 when ps_d1(2) = '1' else    level2 & (3 downto 0 => '0');
   level4 <=  (7 downto 0 => padBit_d1) & level3 when ps_d1(3) = '1' else    level3 & (7 downto 0 => '0');
   level5 <=  (15 downto 0 => padBit_d1) & level4 when ps_d1(4) = '1' else    level4 & (15 downto 0 => '0');
   level6 <=  (31 downto 0 => padBit_d2) & level5_d1 when ps_d2(5) = '1' else    level5_d1 & (31 downto 0 => '0');
   level7 <=  (63 downto 0 => padBit_d2) & level6 when ps_d2(6) = '1' else    level6 & (63 downto 0 => '0');
   level8 <=  (127 downto 0 => padBit_d3) & level7_d1 when ps_d3(7) = '1' else    level7_d1 & (127 downto 0 => '0');
   level9 <=  (255 downto 0 => padBit_d3) & level8 when ps_d3(8) = '1' else    level8 & (255 downto 0 => '0');
   R <= level9(1126 downto 511);
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_1024_F50_uid454
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2016)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: X Y Cin
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_1024_F50_uid454 is
    port (clk : in std_logic;
          X : in  std_logic_vector(1023 downto 0);
          Y : in  std_logic_vector(1023 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(1023 downto 0)   );
end entity;

architecture arch of IntAdder_1024_F50_uid454 is
signal Rtmp :  std_logic_vector(1023 downto 0);
signal Y_d1, Y_d2, Y_d3 :  std_logic_vector(1023 downto 0);
signal Cin_d1, Cin_d2, Cin_d3 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            Y_d1 <=  Y;
            Y_d2 <=  Y_d1;
            Y_d3 <=  Y_d2;
            Cin_d1 <=  Cin;
            Cin_d2 <=  Cin_d1;
            Cin_d3 <=  Cin_d2;
         end if;
      end process;
   Rtmp <= X + Y_d3 + Cin_d3;
   R <= Rtmp;
end architecture;

--------------------------------------------------------------------------------
--                                  PositMAC64
--                    (PositMAC_64_2_Quire_1024_F50_uid2)
-- Inputs: this FMA computes A*B+C
-- VHDL generated for Kintex7 @ 50MHz
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Raul Murillo (2021)
--------------------------------------------------------------------------------
-- Pipeline depth: 3 cycles
-- Clock period (ns): 20
-- Target frequency (MHz): 50
-- Input signals: A B C
-- Output signals: R

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity PositMAC64 is
    port (clk : in std_logic;
          A : in  std_logic_vector(63 downto 0);
          B : in  std_logic_vector(63 downto 0);
          C : in  std_logic_vector(1023 downto 0);
          R : out  std_logic_vector(1023 downto 0)   );
end entity;

architecture arch of PositMAC64 is
   component PositFastDecoder_64_2_F50_uid4 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(63 downto 0);
             Sign : out  std_logic;
             SF : out  std_logic_vector(8 downto 0);
             Frac : out  std_logic_vector(58 downto 0);
             NZN : out  std_logic   );
   end component;

   component PositFastDecoder_64_2_F50_uid8 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(63 downto 0);
             Sign : out  std_logic;
             SF : out  std_logic_vector(8 downto 0);
             Frac : out  std_logic_vector(58 downto 0);
             NZN : out  std_logic   );
   end component;

   component IntMultiplier_F50_uid122 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(60 downto 0);
             Y : in  std_logic_vector(60 downto 0);
             R : out  std_logic_vector(121 downto 0)   );
   end component;

   component IntAdder_10_F50_uid445 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : in  std_logic_vector(9 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(9 downto 0)   );
   end component;

   component IntAdder_10_F50_uid448 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : in  std_logic_vector(9 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(9 downto 0)   );
   end component;

   component IntAdder_9_F50_uid450 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(8 downto 0);
             Y : in  std_logic_vector(8 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(8 downto 0)   );
   end component;

   component RightShifter616_by_max_496_F50_uid452 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(615 downto 0);
             S : in  std_logic_vector(8 downto 0);
             padBit : in  std_logic;
             R : out  std_logic_vector(615 downto 0)   );
   end component;

   component IntAdder_1024_F50_uid454 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(1023 downto 0);
             Y : in  std_logic_vector(1023 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(1023 downto 0)   );
   end component;

signal A_sgn :  std_logic;
signal A_sf :  std_logic_vector(8 downto 0);
signal A_f :  std_logic_vector(58 downto 0);
signal A_nzn :  std_logic;
signal B_sgn :  std_logic;
signal B_sf :  std_logic_vector(8 downto 0);
signal B_f :  std_logic_vector(58 downto 0);
signal B_nzn :  std_logic;
signal AB_nzn, AB_nzn_d1, AB_nzn_d2, AB_nzn_d3 :  std_logic;
signal AB_nar, AB_nar_d1, AB_nar_d2, AB_nar_d3 :  std_logic;
signal AA_f :  std_logic_vector(60 downto 0);
signal BB_f :  std_logic_vector(60 downto 0);
signal AB_f :  std_logic_vector(121 downto 0);
signal AB_sgn, AB_sgn_d1, AB_sgn_d2, AB_sgn_d3 :  std_logic;
signal AB_ovfExtra :  std_logic;
signal AB_ovf :  std_logic;
signal AB_normF :  std_logic_vector(118 downto 0);
signal AA_sf :  std_logic_vector(9 downto 0);
signal BB_sf :  std_logic_vector(9 downto 0);
signal AB_sf_tmp :  std_logic_vector(9 downto 0);
signal AB_sf :  std_logic_vector(9 downto 0);
signal neg_sf, neg_sf_d1, neg_sf_d2, neg_sf_d3 :  std_logic;
signal AB_effectiveSF :  std_logic_vector(8 downto 0);
signal adderInput :  std_logic_vector(8 downto 0);
signal adderBias :  std_logic_vector(8 downto 0);
signal ob :  std_logic;
signal AB_sfBiased :  std_logic_vector(8 downto 0);
signal paddedFrac :  std_logic_vector(615 downto 0);
signal fixedPosit :  std_logic_vector(615 downto 0);
signal quirePosit :  std_logic_vector(992 downto 0);
signal AB_quire :  std_logic_vector(1023 downto 0);
signal zb :  std_logic;
signal ABC_add :  std_logic_vector(1023 downto 0);
signal zeros, zeros_d1, zeros_d2, zeros_d3 :  std_logic_vector(1022 downto 0);
signal C_nar :  std_logic;
signal ABC_nar, ABC_nar_d1, ABC_nar_d2, ABC_nar_d3 :  std_logic;
signal result :  std_logic_vector(1023 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            AB_nzn_d1 <=  AB_nzn;
            AB_nzn_d2 <=  AB_nzn_d1;
            AB_nzn_d3 <=  AB_nzn_d2;
            AB_nar_d1 <=  AB_nar;
            AB_nar_d2 <=  AB_nar_d1;
            AB_nar_d3 <=  AB_nar_d2;
            AB_sgn_d1 <=  AB_sgn;
            AB_sgn_d2 <=  AB_sgn_d1;
            AB_sgn_d3 <=  AB_sgn_d2;
            neg_sf_d1 <=  neg_sf;
            neg_sf_d2 <=  neg_sf_d1;
            neg_sf_d3 <=  neg_sf_d2;
            zeros_d1 <=  zeros;
            zeros_d2 <=  zeros_d1;
            zeros_d3 <=  zeros_d2;
            ABC_nar_d1 <=  ABC_nar;
            ABC_nar_d2 <=  ABC_nar_d1;
            ABC_nar_d3 <=  ABC_nar_d2;
         end if;
      end process;
--------------------------- Start of vhdl generation ---------------------------
---------------------------- Decode A & B operands ----------------------------
   A_decoder: PositFastDecoder_64_2_F50_uid4
      port map ( clk  => clk,
                 X => A,
                 Frac => A_f,
                 NZN => A_nzn,
                 SF => A_sf,
                 Sign => A_sgn);
   B_decoder: PositFastDecoder_64_2_F50_uid8
      port map ( clk  => clk,
                 X => B,
                 Frac => B_f,
                 NZN => B_nzn,
                 SF => B_sf,
                 Sign => B_sgn);
-------------------------------- Multiply A & B --------------------------------
   -- Sign and Special Cases Computation
   AB_nzn <= A_nzn AND B_nzn;
   AB_nar <= (A_sgn AND NOT(A_nzn)) OR (B_sgn AND NOT(B_nzn));
   -- Multiply the fractions
   AA_f <= A_sgn & NOT(A_sgn) & A_f;
   BB_f <= B_sgn & NOT(B_sgn) & B_f;
   FracMultiplier: IntMultiplier_F50_uid122
      port map ( clk  => clk,
                 X => AA_f,
                 Y => BB_f,
                 R => AB_f);
   AB_sgn <= AB_f(121);
   AB_ovfExtra <= NOT(AB_sgn) AND AB_f(120);
   AB_ovf <= AB_ovfExtra OR (AB_sgn XOR AB_f(119));
   AB_normF <= AB_f(118 downto 0) when AB_ovf = '1' else (AB_f(117 downto 0) & '0');
   -- Add the exponent values
   AA_sf <= A_sf(A_sf'high) & A_sf;
   BB_sf <= B_sf(B_sf'high) & B_sf;
   SFAdder: IntAdder_10_F50_uid445
      port map ( clk  => clk,
                 Cin => AB_ovfExtra,
                 X => AA_sf,
                 Y => BB_sf,
                 R => AB_sf_tmp);
   RoundingAdder: IntAdder_10_F50_uid448
      port map ( clk  => clk,
                 Cin => AB_ovf,
                 X => AB_sf_tmp,
                 Y => "0000000000",
                 R => AB_sf);
-------------- Shift AB fraction into corresponding quire format --------------
   neg_sf <= AB_sf(9);
   AB_effectiveSF <= AB_sf(8 downto 0);
   adderInput <= NOT(AB_effectiveSF);
   adderBias <= "111110000" when neg_sf='0' else "111111111";
   ob <= '1';
   BiasedSFAdder: IntAdder_9_F50_uid450
      port map ( clk  => clk,
                 Cin => ob,
                 X => adderInput,
                 Y => adderBias,
                 R => AB_sfBiased);
   paddedFrac <= (NOT(AB_sgn) & AB_normF & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") when neg_sf='0' else ((615 downto 496 => AB_sgn) & NOT(AB_sgn) & AB_normF & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
   Frac_RightShifter: RightShifter616_by_max_496_F50_uid452
      port map ( clk  => clk,
                 S => AB_sfBiased,
                 X => paddedFrac,
                 padBit => AB_sgn,
                 R => fixedPosit);
   quirePosit <= (fixedPosit & "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000") when neg_sf_d3='0' else ((992 downto 616 => AB_sgn_d3) & fixedPosit);
   AB_quire <= ((1023 downto 993 => AB_sgn_d3) & quirePosit) when AB_nzn_d3='1' else AB_nar_d3 & (1022 downto 0 => '0');
---------------------------------- Add quires ----------------------------------
   zb <= '0';
   QuireAdder: IntAdder_1024_F50_uid454
      port map ( clk  => clk,
                 Cin => zb,
                 X => AB_quire,
                 Y => C,
                 R => ABC_add);
   zeros <= (others => '0');
   C_nar <= C(1023) when (C(1022 downto 0) = zeros) else '0';
   ABC_nar <= AB_nar OR C_nar;
   result <= ABC_add when ABC_nar_d3='0' else ('1' & zeros_d3);
   R <= result;
---------------------------- End of vhdl generation ----------------------------
end architecture;

